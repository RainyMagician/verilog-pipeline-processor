
module reg32_0 ( clk, nrst, en, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, nrst, en;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n1;

  DFFX1 \data_out_reg[31]  ( .D(n35), .CLK(clk), .Q(data_out[31]) );
  DFFX1 \data_out_reg[30]  ( .D(n34), .CLK(clk), .Q(data_out[30]) );
  DFFX1 \data_out_reg[29]  ( .D(n33), .CLK(clk), .Q(data_out[29]) );
  DFFX1 \data_out_reg[28]  ( .D(n32), .CLK(clk), .Q(data_out[28]) );
  DFFX1 \data_out_reg[27]  ( .D(n31), .CLK(clk), .Q(data_out[27]) );
  DFFX1 \data_out_reg[26]  ( .D(n30), .CLK(clk), .Q(data_out[26]) );
  DFFX1 \data_out_reg[25]  ( .D(n29), .CLK(clk), .Q(data_out[25]) );
  DFFX1 \data_out_reg[24]  ( .D(n28), .CLK(clk), .Q(data_out[24]) );
  DFFX1 \data_out_reg[23]  ( .D(n27), .CLK(clk), .Q(data_out[23]) );
  DFFX1 \data_out_reg[22]  ( .D(n26), .CLK(clk), .Q(data_out[22]) );
  DFFX1 \data_out_reg[21]  ( .D(n25), .CLK(clk), .Q(data_out[21]) );
  DFFX1 \data_out_reg[20]  ( .D(n24), .CLK(clk), .Q(data_out[20]) );
  DFFX1 \data_out_reg[19]  ( .D(n23), .CLK(clk), .Q(data_out[19]) );
  DFFX1 \data_out_reg[18]  ( .D(n22), .CLK(clk), .Q(data_out[18]) );
  DFFX1 \data_out_reg[17]  ( .D(n21), .CLK(clk), .Q(data_out[17]) );
  DFFX1 \data_out_reg[16]  ( .D(n20), .CLK(clk), .Q(data_out[16]) );
  DFFX1 \data_out_reg[15]  ( .D(n19), .CLK(clk), .Q(data_out[15]) );
  DFFX1 \data_out_reg[14]  ( .D(n18), .CLK(clk), .Q(data_out[14]) );
  DFFX1 \data_out_reg[13]  ( .D(n17), .CLK(clk), .Q(data_out[13]) );
  DFFX1 \data_out_reg[12]  ( .D(n16), .CLK(clk), .Q(data_out[12]) );
  DFFX1 \data_out_reg[11]  ( .D(n15), .CLK(clk), .Q(data_out[11]) );
  DFFX1 \data_out_reg[10]  ( .D(n14), .CLK(clk), .Q(data_out[10]) );
  DFFX1 \data_out_reg[9]  ( .D(n13), .CLK(clk), .Q(data_out[9]) );
  DFFX1 \data_out_reg[8]  ( .D(n12), .CLK(clk), .Q(data_out[8]) );
  DFFX1 \data_out_reg[7]  ( .D(n11), .CLK(clk), .Q(data_out[7]) );
  DFFX1 \data_out_reg[6]  ( .D(n10), .CLK(clk), .Q(data_out[6]) );
  DFFX1 \data_out_reg[5]  ( .D(n9), .CLK(clk), .Q(data_out[5]) );
  DFFX1 \data_out_reg[4]  ( .D(n8), .CLK(clk), .Q(data_out[4]) );
  DFFX1 \data_out_reg[3]  ( .D(n7), .CLK(clk), .Q(data_out[3]) );
  DFFX1 \data_out_reg[2]  ( .D(n6), .CLK(clk), .Q(data_out[2]) );
  DFFX1 \data_out_reg[1]  ( .D(n5), .CLK(clk), .Q(data_out[1]) );
  DFFX1 \data_out_reg[0]  ( .D(n4), .CLK(clk), .Q(data_out[0]) );
  AO22X1 U4 ( .IN1(data_out[0]), .IN2(n2), .IN3(data_in[0]), .IN4(n1), .Q(n4)
         );
  AO22X1 U5 ( .IN1(data_out[1]), .IN2(n2), .IN3(data_in[1]), .IN4(n1), .Q(n5)
         );
  AO22X1 U6 ( .IN1(data_out[2]), .IN2(n2), .IN3(data_in[2]), .IN4(n1), .Q(n6)
         );
  AO22X1 U7 ( .IN1(data_out[3]), .IN2(n2), .IN3(data_in[3]), .IN4(n1), .Q(n7)
         );
  AO22X1 U8 ( .IN1(data_out[4]), .IN2(n2), .IN3(data_in[4]), .IN4(n1), .Q(n8)
         );
  AO22X1 U9 ( .IN1(data_out[5]), .IN2(n2), .IN3(data_in[5]), .IN4(n1), .Q(n9)
         );
  AO22X1 U10 ( .IN1(data_out[6]), .IN2(n2), .IN3(data_in[6]), .IN4(n1), .Q(n10) );
  AO22X1 U11 ( .IN1(data_out[7]), .IN2(n2), .IN3(data_in[7]), .IN4(n1), .Q(n11) );
  AO22X1 U12 ( .IN1(data_out[8]), .IN2(n2), .IN3(data_in[8]), .IN4(n1), .Q(n12) );
  AO22X1 U13 ( .IN1(data_out[9]), .IN2(n2), .IN3(data_in[9]), .IN4(n1), .Q(n13) );
  AO22X1 U14 ( .IN1(data_out[10]), .IN2(n2), .IN3(data_in[10]), .IN4(n1), .Q(
        n14) );
  AO22X1 U15 ( .IN1(data_out[11]), .IN2(n2), .IN3(data_in[11]), .IN4(n1), .Q(
        n15) );
  AO22X1 U16 ( .IN1(data_out[12]), .IN2(n2), .IN3(data_in[12]), .IN4(n1), .Q(
        n16) );
  AO22X1 U17 ( .IN1(data_out[13]), .IN2(n2), .IN3(data_in[13]), .IN4(n1), .Q(
        n17) );
  AO22X1 U18 ( .IN1(data_out[14]), .IN2(n2), .IN3(data_in[14]), .IN4(n1), .Q(
        n18) );
  AO22X1 U19 ( .IN1(data_out[15]), .IN2(n2), .IN3(data_in[15]), .IN4(n1), .Q(
        n19) );
  AO22X1 U20 ( .IN1(data_out[16]), .IN2(n2), .IN3(data_in[16]), .IN4(n1), .Q(
        n20) );
  AO22X1 U21 ( .IN1(data_out[17]), .IN2(n2), .IN3(data_in[17]), .IN4(n1), .Q(
        n21) );
  AO22X1 U22 ( .IN1(data_out[18]), .IN2(n2), .IN3(data_in[18]), .IN4(n1), .Q(
        n22) );
  AO22X1 U23 ( .IN1(data_out[19]), .IN2(n2), .IN3(data_in[19]), .IN4(n1), .Q(
        n23) );
  AO22X1 U24 ( .IN1(data_out[20]), .IN2(n2), .IN3(data_in[20]), .IN4(n1), .Q(
        n24) );
  AO22X1 U25 ( .IN1(data_out[21]), .IN2(n2), .IN3(data_in[21]), .IN4(n1), .Q(
        n25) );
  AO22X1 U26 ( .IN1(data_out[22]), .IN2(n2), .IN3(data_in[22]), .IN4(n1), .Q(
        n26) );
  AO22X1 U27 ( .IN1(data_out[23]), .IN2(n2), .IN3(data_in[23]), .IN4(n1), .Q(
        n27) );
  AO22X1 U28 ( .IN1(data_out[24]), .IN2(n2), .IN3(data_in[24]), .IN4(n1), .Q(
        n28) );
  AO22X1 U29 ( .IN1(data_out[25]), .IN2(n2), .IN3(data_in[25]), .IN4(n1), .Q(
        n29) );
  AO22X1 U30 ( .IN1(data_out[26]), .IN2(n2), .IN3(data_in[26]), .IN4(n1), .Q(
        n30) );
  AO22X1 U31 ( .IN1(data_out[27]), .IN2(n2), .IN3(data_in[27]), .IN4(n1), .Q(
        n31) );
  AO22X1 U32 ( .IN1(data_out[28]), .IN2(n2), .IN3(data_in[28]), .IN4(n1), .Q(
        n32) );
  AO22X1 U33 ( .IN1(data_out[29]), .IN2(n2), .IN3(data_in[29]), .IN4(n1), .Q(
        n33) );
  AO22X1 U34 ( .IN1(data_out[30]), .IN2(n2), .IN3(data_in[30]), .IN4(n1), .Q(
        n34) );
  AO22X1 U35 ( .IN1(data_out[31]), .IN2(n2), .IN3(data_in[31]), .IN4(n1), .Q(
        n35) );
  INVX0 U2 ( .INP(n3), .ZN(n1) );
  AND2X1 U3 ( .IN1(nrst), .IN2(n3), .Q(n2) );
  NAND2X1 U36 ( .IN1(nrst), .IN2(en), .QN(n3) );
endmodule


module if_id_reg ( clk, nrst, en, flush, cur_pc0, next_pc0, cur_pc, next_pc );
  input [31:0] cur_pc0;
  input [31:0] next_pc0;
  output [31:0] cur_pc;
  output [31:0] next_pc;
  input clk, nrst, en, flush;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n1, n2, n69, n70, n71,
         n72, n73;

  DFFX1 \next_pc_reg[31]  ( .D(n68), .CLK(clk), .Q(next_pc[31]) );
  DFFX1 \next_pc_reg[30]  ( .D(n67), .CLK(clk), .Q(next_pc[30]) );
  DFFX1 \next_pc_reg[29]  ( .D(n66), .CLK(clk), .Q(next_pc[29]) );
  DFFX1 \next_pc_reg[28]  ( .D(n65), .CLK(clk), .Q(next_pc[28]) );
  DFFX1 \next_pc_reg[27]  ( .D(n64), .CLK(clk), .Q(next_pc[27]) );
  DFFX1 \next_pc_reg[26]  ( .D(n63), .CLK(clk), .Q(next_pc[26]) );
  DFFX1 \next_pc_reg[25]  ( .D(n62), .CLK(clk), .Q(next_pc[25]) );
  DFFX1 \next_pc_reg[24]  ( .D(n61), .CLK(clk), .Q(next_pc[24]) );
  DFFX1 \next_pc_reg[23]  ( .D(n60), .CLK(clk), .Q(next_pc[23]) );
  DFFX1 \next_pc_reg[22]  ( .D(n59), .CLK(clk), .Q(next_pc[22]) );
  DFFX1 \next_pc_reg[21]  ( .D(n58), .CLK(clk), .Q(next_pc[21]) );
  DFFX1 \next_pc_reg[20]  ( .D(n57), .CLK(clk), .Q(next_pc[20]) );
  DFFX1 \next_pc_reg[19]  ( .D(n56), .CLK(clk), .Q(next_pc[19]) );
  DFFX1 \next_pc_reg[18]  ( .D(n55), .CLK(clk), .Q(next_pc[18]) );
  DFFX1 \next_pc_reg[17]  ( .D(n54), .CLK(clk), .Q(next_pc[17]) );
  DFFX1 \next_pc_reg[16]  ( .D(n53), .CLK(clk), .Q(next_pc[16]) );
  DFFX1 \next_pc_reg[15]  ( .D(n52), .CLK(clk), .Q(next_pc[15]) );
  DFFX1 \next_pc_reg[14]  ( .D(n51), .CLK(clk), .Q(next_pc[14]) );
  DFFX1 \next_pc_reg[13]  ( .D(n50), .CLK(clk), .Q(next_pc[13]) );
  DFFX1 \next_pc_reg[12]  ( .D(n49), .CLK(clk), .Q(next_pc[12]) );
  DFFX1 \next_pc_reg[11]  ( .D(n48), .CLK(clk), .Q(next_pc[11]) );
  DFFX1 \next_pc_reg[10]  ( .D(n47), .CLK(clk), .Q(next_pc[10]) );
  DFFX1 \next_pc_reg[9]  ( .D(n46), .CLK(clk), .Q(next_pc[9]) );
  DFFX1 \next_pc_reg[8]  ( .D(n45), .CLK(clk), .Q(next_pc[8]) );
  DFFX1 \next_pc_reg[7]  ( .D(n44), .CLK(clk), .Q(next_pc[7]) );
  DFFX1 \next_pc_reg[6]  ( .D(n43), .CLK(clk), .Q(next_pc[6]) );
  DFFX1 \next_pc_reg[5]  ( .D(n42), .CLK(clk), .Q(next_pc[5]) );
  DFFX1 \next_pc_reg[4]  ( .D(n41), .CLK(clk), .Q(next_pc[4]) );
  DFFX1 \next_pc_reg[3]  ( .D(n40), .CLK(clk), .Q(next_pc[3]) );
  DFFX1 \next_pc_reg[2]  ( .D(n39), .CLK(clk), .Q(next_pc[2]) );
  DFFX1 \next_pc_reg[1]  ( .D(n38), .CLK(clk), .Q(next_pc[1]) );
  DFFX1 \next_pc_reg[0]  ( .D(n37), .CLK(clk), .Q(next_pc[0]) );
  DFFX1 \cur_pc_reg[31]  ( .D(n36), .CLK(clk), .Q(cur_pc[31]) );
  DFFX1 \cur_pc_reg[30]  ( .D(n35), .CLK(clk), .Q(cur_pc[30]) );
  DFFX1 \cur_pc_reg[29]  ( .D(n34), .CLK(clk), .Q(cur_pc[29]) );
  DFFX1 \cur_pc_reg[28]  ( .D(n33), .CLK(clk), .Q(cur_pc[28]) );
  DFFX1 \cur_pc_reg[27]  ( .D(n32), .CLK(clk), .Q(cur_pc[27]) );
  DFFX1 \cur_pc_reg[26]  ( .D(n31), .CLK(clk), .Q(cur_pc[26]) );
  DFFX1 \cur_pc_reg[25]  ( .D(n30), .CLK(clk), .Q(cur_pc[25]) );
  DFFX1 \cur_pc_reg[24]  ( .D(n29), .CLK(clk), .Q(cur_pc[24]) );
  DFFX1 \cur_pc_reg[23]  ( .D(n28), .CLK(clk), .Q(cur_pc[23]) );
  DFFX1 \cur_pc_reg[22]  ( .D(n27), .CLK(clk), .Q(cur_pc[22]) );
  DFFX1 \cur_pc_reg[21]  ( .D(n26), .CLK(clk), .Q(cur_pc[21]) );
  DFFX1 \cur_pc_reg[20]  ( .D(n25), .CLK(clk), .Q(cur_pc[20]) );
  DFFX1 \cur_pc_reg[19]  ( .D(n24), .CLK(clk), .Q(cur_pc[19]) );
  DFFX1 \cur_pc_reg[18]  ( .D(n23), .CLK(clk), .Q(cur_pc[18]) );
  DFFX1 \cur_pc_reg[17]  ( .D(n22), .CLK(clk), .Q(cur_pc[17]) );
  DFFX1 \cur_pc_reg[16]  ( .D(n21), .CLK(clk), .Q(cur_pc[16]) );
  DFFX1 \cur_pc_reg[15]  ( .D(n20), .CLK(clk), .Q(cur_pc[15]) );
  DFFX1 \cur_pc_reg[14]  ( .D(n19), .CLK(clk), .Q(cur_pc[14]) );
  DFFX1 \cur_pc_reg[13]  ( .D(n18), .CLK(clk), .Q(cur_pc[13]) );
  DFFX1 \cur_pc_reg[12]  ( .D(n17), .CLK(clk), .Q(cur_pc[12]) );
  DFFX1 \cur_pc_reg[11]  ( .D(n16), .CLK(clk), .Q(cur_pc[11]) );
  DFFX1 \cur_pc_reg[10]  ( .D(n15), .CLK(clk), .Q(cur_pc[10]) );
  DFFX1 \cur_pc_reg[9]  ( .D(n14), .CLK(clk), .Q(cur_pc[9]) );
  DFFX1 \cur_pc_reg[8]  ( .D(n13), .CLK(clk), .Q(cur_pc[8]) );
  DFFX1 \cur_pc_reg[7]  ( .D(n12), .CLK(clk), .Q(cur_pc[7]) );
  DFFX1 \cur_pc_reg[6]  ( .D(n11), .CLK(clk), .Q(cur_pc[6]) );
  DFFX1 \cur_pc_reg[5]  ( .D(n10), .CLK(clk), .Q(cur_pc[5]) );
  DFFX1 \cur_pc_reg[4]  ( .D(n9), .CLK(clk), .Q(cur_pc[4]) );
  DFFX1 \cur_pc_reg[3]  ( .D(n8), .CLK(clk), .Q(cur_pc[3]) );
  DFFX1 \cur_pc_reg[2]  ( .D(n7), .CLK(clk), .Q(cur_pc[2]) );
  DFFX1 \cur_pc_reg[1]  ( .D(n6), .CLK(clk), .Q(cur_pc[1]) );
  DFFX1 \cur_pc_reg[0]  ( .D(n5), .CLK(clk), .Q(cur_pc[0]) );
  AO22X1 U4 ( .IN1(cur_pc[0]), .IN2(n3), .IN3(cur_pc0[0]), .IN4(n72), .Q(n5)
         );
  AO22X1 U5 ( .IN1(cur_pc[1]), .IN2(n3), .IN3(cur_pc0[1]), .IN4(n72), .Q(n6)
         );
  AO22X1 U6 ( .IN1(cur_pc[2]), .IN2(n3), .IN3(cur_pc0[2]), .IN4(n72), .Q(n7)
         );
  AO22X1 U7 ( .IN1(cur_pc[3]), .IN2(n3), .IN3(cur_pc0[3]), .IN4(n72), .Q(n8)
         );
  AO22X1 U8 ( .IN1(cur_pc[4]), .IN2(n3), .IN3(cur_pc0[4]), .IN4(n72), .Q(n9)
         );
  AO22X1 U9 ( .IN1(cur_pc[5]), .IN2(n3), .IN3(cur_pc0[5]), .IN4(n72), .Q(n10)
         );
  AO22X1 U10 ( .IN1(cur_pc[6]), .IN2(n3), .IN3(cur_pc0[6]), .IN4(n72), .Q(n11)
         );
  AO22X1 U11 ( .IN1(cur_pc[7]), .IN2(n3), .IN3(cur_pc0[7]), .IN4(n72), .Q(n12)
         );
  AO22X1 U12 ( .IN1(cur_pc[8]), .IN2(n3), .IN3(cur_pc0[8]), .IN4(n72), .Q(n13)
         );
  AO22X1 U13 ( .IN1(cur_pc[9]), .IN2(n3), .IN3(cur_pc0[9]), .IN4(n72), .Q(n14)
         );
  AO22X1 U14 ( .IN1(cur_pc[10]), .IN2(n3), .IN3(cur_pc0[10]), .IN4(n72), .Q(
        n15) );
  AO22X1 U15 ( .IN1(cur_pc[11]), .IN2(n3), .IN3(cur_pc0[11]), .IN4(n72), .Q(
        n16) );
  AO22X1 U16 ( .IN1(cur_pc[12]), .IN2(n1), .IN3(cur_pc0[12]), .IN4(n72), .Q(
        n17) );
  AO22X1 U17 ( .IN1(cur_pc[13]), .IN2(n1), .IN3(cur_pc0[13]), .IN4(n72), .Q(
        n18) );
  AO22X1 U18 ( .IN1(cur_pc[14]), .IN2(n1), .IN3(cur_pc0[14]), .IN4(n72), .Q(
        n19) );
  AO22X1 U19 ( .IN1(cur_pc[15]), .IN2(n1), .IN3(cur_pc0[15]), .IN4(n72), .Q(
        n20) );
  AO22X1 U20 ( .IN1(cur_pc[16]), .IN2(n1), .IN3(cur_pc0[16]), .IN4(n72), .Q(
        n21) );
  AO22X1 U21 ( .IN1(cur_pc[17]), .IN2(n1), .IN3(cur_pc0[17]), .IN4(n72), .Q(
        n22) );
  AO22X1 U22 ( .IN1(cur_pc[18]), .IN2(n1), .IN3(cur_pc0[18]), .IN4(n72), .Q(
        n23) );
  AO22X1 U23 ( .IN1(cur_pc[19]), .IN2(n1), .IN3(cur_pc0[19]), .IN4(n72), .Q(
        n24) );
  AO22X1 U24 ( .IN1(cur_pc[20]), .IN2(n1), .IN3(cur_pc0[20]), .IN4(n72), .Q(
        n25) );
  AO22X1 U25 ( .IN1(cur_pc[21]), .IN2(n1), .IN3(cur_pc0[21]), .IN4(n72), .Q(
        n26) );
  AO22X1 U26 ( .IN1(cur_pc[22]), .IN2(n1), .IN3(cur_pc0[22]), .IN4(n72), .Q(
        n27) );
  AO22X1 U27 ( .IN1(cur_pc[23]), .IN2(n1), .IN3(cur_pc0[23]), .IN4(n72), .Q(
        n28) );
  AO22X1 U28 ( .IN1(cur_pc[24]), .IN2(n2), .IN3(cur_pc0[24]), .IN4(n72), .Q(
        n29) );
  AO22X1 U29 ( .IN1(cur_pc[25]), .IN2(n2), .IN3(cur_pc0[25]), .IN4(n72), .Q(
        n30) );
  AO22X1 U30 ( .IN1(cur_pc[26]), .IN2(n2), .IN3(cur_pc0[26]), .IN4(n72), .Q(
        n31) );
  AO22X1 U31 ( .IN1(cur_pc[27]), .IN2(n2), .IN3(cur_pc0[27]), .IN4(n72), .Q(
        n32) );
  AO22X1 U32 ( .IN1(cur_pc[28]), .IN2(n2), .IN3(cur_pc0[28]), .IN4(n72), .Q(
        n33) );
  AO22X1 U33 ( .IN1(cur_pc[29]), .IN2(n2), .IN3(cur_pc0[29]), .IN4(n72), .Q(
        n34) );
  AO22X1 U34 ( .IN1(cur_pc[30]), .IN2(n2), .IN3(cur_pc0[30]), .IN4(n72), .Q(
        n35) );
  AO22X1 U35 ( .IN1(cur_pc[31]), .IN2(n2), .IN3(cur_pc0[31]), .IN4(n72), .Q(
        n36) );
  AO22X1 U36 ( .IN1(next_pc[0]), .IN2(n2), .IN3(next_pc0[0]), .IN4(n72), .Q(
        n37) );
  AO22X1 U37 ( .IN1(next_pc[1]), .IN2(n2), .IN3(next_pc0[1]), .IN4(n72), .Q(
        n38) );
  AO22X1 U38 ( .IN1(next_pc[2]), .IN2(n2), .IN3(next_pc0[2]), .IN4(n72), .Q(
        n39) );
  AO22X1 U39 ( .IN1(next_pc[3]), .IN2(n2), .IN3(next_pc0[3]), .IN4(n72), .Q(
        n40) );
  AO22X1 U40 ( .IN1(next_pc[4]), .IN2(n69), .IN3(next_pc0[4]), .IN4(n72), .Q(
        n41) );
  AO22X1 U41 ( .IN1(next_pc[5]), .IN2(n69), .IN3(next_pc0[5]), .IN4(n72), .Q(
        n42) );
  AO22X1 U42 ( .IN1(next_pc[6]), .IN2(n69), .IN3(next_pc0[6]), .IN4(n72), .Q(
        n43) );
  AO22X1 U43 ( .IN1(next_pc[7]), .IN2(n69), .IN3(next_pc0[7]), .IN4(n72), .Q(
        n44) );
  AO22X1 U44 ( .IN1(next_pc[8]), .IN2(n69), .IN3(next_pc0[8]), .IN4(n72), .Q(
        n45) );
  AO22X1 U45 ( .IN1(next_pc[9]), .IN2(n69), .IN3(next_pc0[9]), .IN4(n72), .Q(
        n46) );
  AO22X1 U46 ( .IN1(next_pc[10]), .IN2(n69), .IN3(next_pc0[10]), .IN4(n72), 
        .Q(n47) );
  AO22X1 U47 ( .IN1(next_pc[11]), .IN2(n69), .IN3(next_pc0[11]), .IN4(n72), 
        .Q(n48) );
  AO22X1 U48 ( .IN1(next_pc[12]), .IN2(n69), .IN3(next_pc0[12]), .IN4(n72), 
        .Q(n49) );
  AO22X1 U49 ( .IN1(next_pc[13]), .IN2(n69), .IN3(next_pc0[13]), .IN4(n72), 
        .Q(n50) );
  AO22X1 U50 ( .IN1(next_pc[14]), .IN2(n69), .IN3(next_pc0[14]), .IN4(n72), 
        .Q(n51) );
  AO22X1 U51 ( .IN1(next_pc[15]), .IN2(n69), .IN3(next_pc0[15]), .IN4(n72), 
        .Q(n52) );
  AO22X1 U52 ( .IN1(next_pc[16]), .IN2(n70), .IN3(next_pc0[16]), .IN4(n72), 
        .Q(n53) );
  AO22X1 U53 ( .IN1(next_pc[17]), .IN2(n70), .IN3(next_pc0[17]), .IN4(n72), 
        .Q(n54) );
  AO22X1 U54 ( .IN1(next_pc[18]), .IN2(n70), .IN3(next_pc0[18]), .IN4(n72), 
        .Q(n55) );
  AO22X1 U55 ( .IN1(next_pc[19]), .IN2(n70), .IN3(next_pc0[19]), .IN4(n72), 
        .Q(n56) );
  AO22X1 U56 ( .IN1(next_pc[20]), .IN2(n70), .IN3(next_pc0[20]), .IN4(n72), 
        .Q(n57) );
  AO22X1 U57 ( .IN1(next_pc[21]), .IN2(n70), .IN3(next_pc0[21]), .IN4(n72), 
        .Q(n58) );
  AO22X1 U58 ( .IN1(next_pc[22]), .IN2(n70), .IN3(next_pc0[22]), .IN4(n72), 
        .Q(n59) );
  AO22X1 U59 ( .IN1(next_pc[23]), .IN2(n70), .IN3(next_pc0[23]), .IN4(n72), 
        .Q(n60) );
  AO22X1 U60 ( .IN1(next_pc[24]), .IN2(n70), .IN3(next_pc0[24]), .IN4(n72), 
        .Q(n61) );
  AO22X1 U61 ( .IN1(next_pc[25]), .IN2(n70), .IN3(next_pc0[25]), .IN4(n72), 
        .Q(n62) );
  AO22X1 U62 ( .IN1(next_pc[26]), .IN2(n70), .IN3(next_pc0[26]), .IN4(n72), 
        .Q(n63) );
  AO22X1 U63 ( .IN1(next_pc[27]), .IN2(n70), .IN3(next_pc0[27]), .IN4(n72), 
        .Q(n64) );
  AO22X1 U64 ( .IN1(next_pc[28]), .IN2(n3), .IN3(next_pc0[28]), .IN4(n72), .Q(
        n65) );
  AO22X1 U65 ( .IN1(next_pc[29]), .IN2(n3), .IN3(next_pc0[29]), .IN4(n72), .Q(
        n66) );
  AO22X1 U66 ( .IN1(next_pc[30]), .IN2(n3), .IN3(next_pc0[30]), .IN4(n72), .Q(
        n67) );
  AO22X1 U67 ( .IN1(next_pc[31]), .IN2(n3), .IN3(next_pc0[31]), .IN4(n72), .Q(
        n68) );
  AND3X1 U68 ( .IN1(n4), .IN2(n73), .IN3(nrst), .Q(n3) );
  NAND3X0 U69 ( .IN1(en), .IN2(n73), .IN3(nrst), .QN(n4) );
  INVX0 U2 ( .INP(n3), .ZN(n71) );
  INVX0 U3 ( .INP(flush), .ZN(n73) );
  INVX0 U70 ( .INP(n71), .ZN(n1) );
  INVX0 U71 ( .INP(n71), .ZN(n2) );
  INVX0 U72 ( .INP(n71), .ZN(n69) );
  INVX0 U73 ( .INP(n71), .ZN(n70) );
  INVX2 U74 ( .INP(n4), .ZN(n72) );
endmodule


module rf ( clk, nrst, wr_en, rd_addrA, rd_addrB, wr_addr, wr_data, rd_dataA, 
        rd_dataB );
  input [4:0] rd_addrA;
  input [4:0] rd_addrB;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_dataA;
  output [31:0] rd_dataB;
  input clk, nrst, wr_en;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, \mem[31][31] ,
         \mem[31][30] , \mem[31][29] , \mem[31][28] , \mem[31][27] ,
         \mem[31][26] , \mem[31][25] , \mem[31][24] , \mem[31][23] ,
         \mem[31][22] , \mem[31][21] , \mem[31][20] , \mem[31][19] ,
         \mem[31][18] , \mem[31][17] , \mem[31][16] , \mem[31][15] ,
         \mem[31][14] , \mem[31][13] , \mem[31][12] , \mem[31][11] ,
         \mem[31][10] , \mem[31][9] , \mem[31][8] , \mem[31][7] , \mem[31][6] ,
         \mem[31][5] , \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] ,
         \mem[31][0] , \mem[30][31] , \mem[30][30] , \mem[30][29] ,
         \mem[30][28] , \mem[30][27] , \mem[30][26] , \mem[30][25] ,
         \mem[30][24] , \mem[30][23] , \mem[30][22] , \mem[30][21] ,
         \mem[30][20] , \mem[30][19] , \mem[30][18] , \mem[30][17] ,
         \mem[30][16] , \mem[30][15] , \mem[30][14] , \mem[30][13] ,
         \mem[30][12] , \mem[30][11] , \mem[30][10] , \mem[30][9] ,
         \mem[30][8] , \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] ,
         \mem[30][3] , \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][31] ,
         \mem[29][30] , \mem[29][29] , \mem[29][28] , \mem[29][27] ,
         \mem[29][26] , \mem[29][25] , \mem[29][24] , \mem[29][23] ,
         \mem[29][22] , \mem[29][21] , \mem[29][20] , \mem[29][19] ,
         \mem[29][18] , \mem[29][17] , \mem[29][16] , \mem[29][15] ,
         \mem[29][14] , \mem[29][13] , \mem[29][12] , \mem[29][11] ,
         \mem[29][10] , \mem[29][9] , \mem[29][8] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][31] , \mem[28][30] , \mem[28][29] ,
         \mem[28][28] , \mem[28][27] , \mem[28][26] , \mem[28][25] ,
         \mem[28][24] , \mem[28][23] , \mem[28][22] , \mem[28][21] ,
         \mem[28][20] , \mem[28][19] , \mem[28][18] , \mem[28][17] ,
         \mem[28][16] , \mem[28][15] , \mem[28][14] , \mem[28][13] ,
         \mem[28][12] , \mem[28][11] , \mem[28][10] , \mem[28][9] ,
         \mem[28][8] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][31] ,
         \mem[27][30] , \mem[27][29] , \mem[27][28] , \mem[27][27] ,
         \mem[27][26] , \mem[27][25] , \mem[27][24] , \mem[27][23] ,
         \mem[27][22] , \mem[27][21] , \mem[27][20] , \mem[27][19] ,
         \mem[27][18] , \mem[27][17] , \mem[27][16] , \mem[27][15] ,
         \mem[27][14] , \mem[27][13] , \mem[27][12] , \mem[27][11] ,
         \mem[27][10] , \mem[27][9] , \mem[27][8] , \mem[27][7] , \mem[27][6] ,
         \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] , \mem[27][1] ,
         \mem[27][0] , \mem[26][31] , \mem[26][30] , \mem[26][29] ,
         \mem[26][28] , \mem[26][27] , \mem[26][26] , \mem[26][25] ,
         \mem[26][24] , \mem[26][23] , \mem[26][22] , \mem[26][21] ,
         \mem[26][20] , \mem[26][19] , \mem[26][18] , \mem[26][17] ,
         \mem[26][16] , \mem[26][15] , \mem[26][14] , \mem[26][13] ,
         \mem[26][12] , \mem[26][11] , \mem[26][10] , \mem[26][9] ,
         \mem[26][8] , \mem[26][7] , \mem[26][6] , \mem[26][5] , \mem[26][4] ,
         \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] , \mem[25][31] ,
         \mem[25][30] , \mem[25][29] , \mem[25][28] , \mem[25][27] ,
         \mem[25][26] , \mem[25][25] , \mem[25][24] , \mem[25][23] ,
         \mem[25][22] , \mem[25][21] , \mem[25][20] , \mem[25][19] ,
         \mem[25][18] , \mem[25][17] , \mem[25][16] , \mem[25][15] ,
         \mem[25][14] , \mem[25][13] , \mem[25][12] , \mem[25][11] ,
         \mem[25][10] , \mem[25][9] , \mem[25][8] , \mem[25][7] , \mem[25][6] ,
         \mem[25][5] , \mem[25][4] , \mem[25][3] , \mem[25][2] , \mem[25][1] ,
         \mem[25][0] , \mem[24][31] , \mem[24][30] , \mem[24][29] ,
         \mem[24][28] , \mem[24][27] , \mem[24][26] , \mem[24][25] ,
         \mem[24][24] , \mem[24][23] , \mem[24][22] , \mem[24][21] ,
         \mem[24][20] , \mem[24][19] , \mem[24][18] , \mem[24][17] ,
         \mem[24][16] , \mem[24][15] , \mem[24][14] , \mem[24][13] ,
         \mem[24][12] , \mem[24][11] , \mem[24][10] , \mem[24][9] ,
         \mem[24][8] , \mem[24][7] , \mem[24][6] , \mem[24][5] , \mem[24][4] ,
         \mem[24][3] , \mem[24][2] , \mem[24][1] , \mem[24][0] , \mem[23][31] ,
         \mem[23][30] , \mem[23][29] , \mem[23][28] , \mem[23][27] ,
         \mem[23][26] , \mem[23][25] , \mem[23][24] , \mem[23][23] ,
         \mem[23][22] , \mem[23][21] , \mem[23][20] , \mem[23][19] ,
         \mem[23][18] , \mem[23][17] , \mem[23][16] , \mem[23][15] ,
         \mem[23][14] , \mem[23][13] , \mem[23][12] , \mem[23][11] ,
         \mem[23][10] , \mem[23][9] , \mem[23][8] , \mem[23][7] , \mem[23][6] ,
         \mem[23][5] , \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] ,
         \mem[23][0] , \mem[22][31] , \mem[22][30] , \mem[22][29] ,
         \mem[22][28] , \mem[22][27] , \mem[22][26] , \mem[22][25] ,
         \mem[22][24] , \mem[22][23] , \mem[22][22] , \mem[22][21] ,
         \mem[22][20] , \mem[22][19] , \mem[22][18] , \mem[22][17] ,
         \mem[22][16] , \mem[22][15] , \mem[22][14] , \mem[22][13] ,
         \mem[22][12] , \mem[22][11] , \mem[22][10] , \mem[22][9] ,
         \mem[22][8] , \mem[22][7] , \mem[22][6] , \mem[22][5] , \mem[22][4] ,
         \mem[22][3] , \mem[22][2] , \mem[22][1] , \mem[22][0] , \mem[21][31] ,
         \mem[21][30] , \mem[21][29] , \mem[21][28] , \mem[21][27] ,
         \mem[21][26] , \mem[21][25] , \mem[21][24] , \mem[21][23] ,
         \mem[21][22] , \mem[21][21] , \mem[21][20] , \mem[21][19] ,
         \mem[21][18] , \mem[21][17] , \mem[21][16] , \mem[21][15] ,
         \mem[21][14] , \mem[21][13] , \mem[21][12] , \mem[21][11] ,
         \mem[21][10] , \mem[21][9] , \mem[21][8] , \mem[21][7] , \mem[21][6] ,
         \mem[21][5] , \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] ,
         \mem[21][0] , \mem[20][31] , \mem[20][30] , \mem[20][29] ,
         \mem[20][28] , \mem[20][27] , \mem[20][26] , \mem[20][25] ,
         \mem[20][24] , \mem[20][23] , \mem[20][22] , \mem[20][21] ,
         \mem[20][20] , \mem[20][19] , \mem[20][18] , \mem[20][17] ,
         \mem[20][16] , \mem[20][15] , \mem[20][14] , \mem[20][13] ,
         \mem[20][12] , \mem[20][11] , \mem[20][10] , \mem[20][9] ,
         \mem[20][8] , \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] ,
         \mem[20][3] , \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][31] ,
         \mem[19][30] , \mem[19][29] , \mem[19][28] , \mem[19][27] ,
         \mem[19][26] , \mem[19][25] , \mem[19][24] , \mem[19][23] ,
         \mem[19][22] , \mem[19][21] , \mem[19][20] , \mem[19][19] ,
         \mem[19][18] , \mem[19][17] , \mem[19][16] , \mem[19][15] ,
         \mem[19][14] , \mem[19][13] , \mem[19][12] , \mem[19][11] ,
         \mem[19][10] , \mem[19][9] , \mem[19][8] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][31] , \mem[18][30] , \mem[18][29] ,
         \mem[18][28] , \mem[18][27] , \mem[18][26] , \mem[18][25] ,
         \mem[18][24] , \mem[18][23] , \mem[18][22] , \mem[18][21] ,
         \mem[18][20] , \mem[18][19] , \mem[18][18] , \mem[18][17] ,
         \mem[18][16] , \mem[18][15] , \mem[18][14] , \mem[18][13] ,
         \mem[18][12] , \mem[18][11] , \mem[18][10] , \mem[18][9] ,
         \mem[18][8] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][31] ,
         \mem[17][30] , \mem[17][29] , \mem[17][28] , \mem[17][27] ,
         \mem[17][26] , \mem[17][25] , \mem[17][24] , \mem[17][23] ,
         \mem[17][22] , \mem[17][21] , \mem[17][20] , \mem[17][19] ,
         \mem[17][18] , \mem[17][17] , \mem[17][16] , \mem[17][15] ,
         \mem[17][14] , \mem[17][13] , \mem[17][12] , \mem[17][11] ,
         \mem[17][10] , \mem[17][9] , \mem[17][8] , \mem[17][7] , \mem[17][6] ,
         \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] , \mem[17][1] ,
         \mem[17][0] , \mem[16][31] , \mem[16][30] , \mem[16][29] ,
         \mem[16][28] , \mem[16][27] , \mem[16][26] , \mem[16][25] ,
         \mem[16][24] , \mem[16][23] , \mem[16][22] , \mem[16][21] ,
         \mem[16][20] , \mem[16][19] , \mem[16][18] , \mem[16][17] ,
         \mem[16][16] , \mem[16][15] , \mem[16][14] , \mem[16][13] ,
         \mem[16][12] , \mem[16][11] , \mem[16][10] , \mem[16][9] ,
         \mem[16][8] , \mem[16][7] , \mem[16][6] , \mem[16][5] , \mem[16][4] ,
         \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] , \mem[15][31] ,
         \mem[15][30] , \mem[15][29] , \mem[15][28] , \mem[15][27] ,
         \mem[15][26] , \mem[15][25] , \mem[15][24] , \mem[15][23] ,
         \mem[15][22] , \mem[15][21] , \mem[15][20] , \mem[15][19] ,
         \mem[15][18] , \mem[15][17] , \mem[15][16] , \mem[15][15] ,
         \mem[15][14] , \mem[15][13] , \mem[15][12] , \mem[15][11] ,
         \mem[15][10] , \mem[15][9] , \mem[15][8] , \mem[15][7] , \mem[15][6] ,
         \mem[15][5] , \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] ,
         \mem[15][0] , \mem[14][31] , \mem[14][30] , \mem[14][29] ,
         \mem[14][28] , \mem[14][27] , \mem[14][26] , \mem[14][25] ,
         \mem[14][24] , \mem[14][23] , \mem[14][22] , \mem[14][21] ,
         \mem[14][20] , \mem[14][19] , \mem[14][18] , \mem[14][17] ,
         \mem[14][16] , \mem[14][15] , \mem[14][14] , \mem[14][13] ,
         \mem[14][12] , \mem[14][11] , \mem[14][10] , \mem[14][9] ,
         \mem[14][8] , \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] ,
         \mem[14][3] , \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][31] ,
         \mem[13][30] , \mem[13][29] , \mem[13][28] , \mem[13][27] ,
         \mem[13][26] , \mem[13][25] , \mem[13][24] , \mem[13][23] ,
         \mem[13][22] , \mem[13][21] , \mem[13][20] , \mem[13][19] ,
         \mem[13][18] , \mem[13][17] , \mem[13][16] , \mem[13][15] ,
         \mem[13][14] , \mem[13][13] , \mem[13][12] , \mem[13][11] ,
         \mem[13][10] , \mem[13][9] , \mem[13][8] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][31] , \mem[12][30] , \mem[12][29] ,
         \mem[12][28] , \mem[12][27] , \mem[12][26] , \mem[12][25] ,
         \mem[12][24] , \mem[12][23] , \mem[12][22] , \mem[12][21] ,
         \mem[12][20] , \mem[12][19] , \mem[12][18] , \mem[12][17] ,
         \mem[12][16] , \mem[12][15] , \mem[12][14] , \mem[12][13] ,
         \mem[12][12] , \mem[12][11] , \mem[12][10] , \mem[12][9] ,
         \mem[12][8] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][31] ,
         \mem[11][30] , \mem[11][29] , \mem[11][28] , \mem[11][27] ,
         \mem[11][26] , \mem[11][25] , \mem[11][24] , \mem[11][23] ,
         \mem[11][22] , \mem[11][21] , \mem[11][20] , \mem[11][19] ,
         \mem[11][18] , \mem[11][17] , \mem[11][16] , \mem[11][15] ,
         \mem[11][14] , \mem[11][13] , \mem[11][12] , \mem[11][11] ,
         \mem[11][10] , \mem[11][9] , \mem[11][8] , \mem[11][7] , \mem[11][6] ,
         \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] ,
         \mem[11][0] , \mem[10][31] , \mem[10][30] , \mem[10][29] ,
         \mem[10][28] , \mem[10][27] , \mem[10][26] , \mem[10][25] ,
         \mem[10][24] , \mem[10][23] , \mem[10][22] , \mem[10][21] ,
         \mem[10][20] , \mem[10][19] , \mem[10][18] , \mem[10][17] ,
         \mem[10][16] , \mem[10][15] , \mem[10][14] , \mem[10][13] ,
         \mem[10][12] , \mem[10][11] , \mem[10][10] , \mem[10][9] ,
         \mem[10][8] , \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] ,
         \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][31] ,
         \mem[9][30] , \mem[9][29] , \mem[9][28] , \mem[9][27] , \mem[9][26] ,
         \mem[9][25] , \mem[9][24] , \mem[9][23] , \mem[9][22] , \mem[9][21] ,
         \mem[9][20] , \mem[9][19] , \mem[9][18] , \mem[9][17] , \mem[9][16] ,
         \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] , \mem[9][11] ,
         \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][31] , \mem[8][30] , \mem[8][29] , \mem[8][28] ,
         \mem[8][27] , \mem[8][26] , \mem[8][25] , \mem[8][24] , \mem[8][23] ,
         \mem[8][22] , \mem[8][21] , \mem[8][20] , \mem[8][19] , \mem[8][18] ,
         \mem[8][17] , \mem[8][16] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][31] , \mem[7][30] ,
         \mem[7][29] , \mem[7][28] , \mem[7][27] , \mem[7][26] , \mem[7][25] ,
         \mem[7][24] , \mem[7][23] , \mem[7][22] , \mem[7][21] , \mem[7][20] ,
         \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] , \mem[7][15] ,
         \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] ,
         \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] ,
         \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] ,
         \mem[6][31] , \mem[6][30] , \mem[6][29] , \mem[6][28] , \mem[6][27] ,
         \mem[6][26] , \mem[6][25] , \mem[6][24] , \mem[6][23] , \mem[6][22] ,
         \mem[6][21] , \mem[6][20] , \mem[6][19] , \mem[6][18] , \mem[6][17] ,
         \mem[6][16] , \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] ,
         \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][31] , \mem[5][30] , \mem[5][29] ,
         \mem[5][28] , \mem[5][27] , \mem[5][26] , \mem[5][25] , \mem[5][24] ,
         \mem[5][23] , \mem[5][22] , \mem[5][21] , \mem[5][20] , \mem[5][19] ,
         \mem[5][18] , \mem[5][17] , \mem[5][16] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][31] ,
         \mem[4][30] , \mem[4][29] , \mem[4][28] , \mem[4][27] , \mem[4][26] ,
         \mem[4][25] , \mem[4][24] , \mem[4][23] , \mem[4][22] , \mem[4][21] ,
         \mem[4][20] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][31] , \mem[3][30] , \mem[3][29] , \mem[3][28] ,
         \mem[3][27] , \mem[3][26] , \mem[3][25] , \mem[3][24] , \mem[3][23] ,
         \mem[3][22] , \mem[3][21] , \mem[3][20] , \mem[3][19] , \mem[3][18] ,
         \mem[3][17] , \mem[3][16] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][31] , \mem[2][30] ,
         \mem[2][29] , \mem[2][28] , \mem[2][27] , \mem[2][26] , \mem[2][25] ,
         \mem[2][24] , \mem[2][23] , \mem[2][22] , \mem[2][21] , \mem[2][20] ,
         \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] , \mem[2][15] ,
         \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] ,
         \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] ,
         \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] ,
         \mem[1][31] , \mem[1][30] , \mem[1][29] , \mem[1][28] , \mem[1][27] ,
         \mem[1][26] , \mem[1][25] , \mem[1][24] , \mem[1][23] , \mem[1][22] ,
         \mem[1][21] , \mem[1][20] , \mem[1][19] , \mem[1][18] , \mem[1][17] ,
         \mem[1][16] , \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] ,
         \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][31] , \mem[0][30] , \mem[0][29] ,
         \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] , \mem[0][24] ,
         \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] ,
         \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n92, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004;
  assign N10 = rd_addrA[0];
  assign N11 = rd_addrA[1];
  assign N12 = rd_addrA[2];
  assign N13 = rd_addrA[3];
  assign N14 = rd_addrA[4];
  assign N15 = rd_addrB[0];
  assign N16 = rd_addrB[1];
  assign N17 = rd_addrB[2];
  assign N18 = rd_addrB[3];
  assign N19 = rd_addrB[4];

  DFFX1 \mem_reg[31][31]  ( .D(n1137), .CLK(clk), .Q(\mem[31][31] ) );
  DFFX1 \mem_reg[31][30]  ( .D(n1136), .CLK(clk), .Q(\mem[31][30] ) );
  DFFX1 \mem_reg[31][29]  ( .D(n1135), .CLK(clk), .Q(\mem[31][29] ) );
  DFFX1 \mem_reg[31][28]  ( .D(n1134), .CLK(clk), .Q(\mem[31][28] ) );
  DFFX1 \mem_reg[31][27]  ( .D(n1133), .CLK(clk), .Q(\mem[31][27] ) );
  DFFX1 \mem_reg[31][26]  ( .D(n1132), .CLK(clk), .Q(\mem[31][26] ) );
  DFFX1 \mem_reg[31][25]  ( .D(n1131), .CLK(clk), .Q(\mem[31][25] ) );
  DFFX1 \mem_reg[31][24]  ( .D(n1130), .CLK(clk), .Q(\mem[31][24] ) );
  DFFX1 \mem_reg[31][23]  ( .D(n1129), .CLK(clk), .Q(\mem[31][23] ) );
  DFFX1 \mem_reg[31][22]  ( .D(n1128), .CLK(clk), .Q(\mem[31][22] ) );
  DFFX1 \mem_reg[31][21]  ( .D(n1127), .CLK(clk), .Q(\mem[31][21] ) );
  DFFX1 \mem_reg[31][20]  ( .D(n1126), .CLK(clk), .Q(\mem[31][20] ) );
  DFFX1 \mem_reg[31][19]  ( .D(n1125), .CLK(clk), .Q(\mem[31][19] ) );
  DFFX1 \mem_reg[31][18]  ( .D(n1124), .CLK(clk), .Q(\mem[31][18] ) );
  DFFX1 \mem_reg[31][17]  ( .D(n1123), .CLK(clk), .Q(\mem[31][17] ) );
  DFFX1 \mem_reg[31][16]  ( .D(n1122), .CLK(clk), .Q(\mem[31][16] ) );
  DFFX1 \mem_reg[31][15]  ( .D(n1121), .CLK(clk), .Q(\mem[31][15] ) );
  DFFX1 \mem_reg[31][14]  ( .D(n1120), .CLK(clk), .Q(\mem[31][14] ) );
  DFFX1 \mem_reg[31][13]  ( .D(n1119), .CLK(clk), .Q(\mem[31][13] ) );
  DFFX1 \mem_reg[31][12]  ( .D(n1118), .CLK(clk), .Q(\mem[31][12] ) );
  DFFX1 \mem_reg[31][11]  ( .D(n1117), .CLK(clk), .Q(\mem[31][11] ) );
  DFFX1 \mem_reg[31][10]  ( .D(n1116), .CLK(clk), .Q(\mem[31][10] ) );
  DFFX1 \mem_reg[31][9]  ( .D(n1115), .CLK(clk), .Q(\mem[31][9] ) );
  DFFX1 \mem_reg[31][8]  ( .D(n1114), .CLK(clk), .Q(\mem[31][8] ) );
  DFFX1 \mem_reg[31][7]  ( .D(n1113), .CLK(clk), .Q(\mem[31][7] ) );
  DFFX1 \mem_reg[31][6]  ( .D(n1112), .CLK(clk), .Q(\mem[31][6] ) );
  DFFX1 \mem_reg[31][5]  ( .D(n1111), .CLK(clk), .Q(\mem[31][5] ) );
  DFFX1 \mem_reg[31][4]  ( .D(n1110), .CLK(clk), .Q(\mem[31][4] ) );
  DFFX1 \mem_reg[31][3]  ( .D(n1109), .CLK(clk), .Q(\mem[31][3] ) );
  DFFX1 \mem_reg[31][2]  ( .D(n1108), .CLK(clk), .Q(\mem[31][2] ) );
  DFFX1 \mem_reg[31][1]  ( .D(n1107), .CLK(clk), .Q(\mem[31][1] ) );
  DFFX1 \mem_reg[31][0]  ( .D(n1106), .CLK(clk), .Q(\mem[31][0] ) );
  DFFX1 \mem_reg[30][31]  ( .D(n1105), .CLK(clk), .Q(\mem[30][31] ) );
  DFFX1 \mem_reg[30][30]  ( .D(n1104), .CLK(clk), .Q(\mem[30][30] ) );
  DFFX1 \mem_reg[30][29]  ( .D(n1103), .CLK(clk), .Q(\mem[30][29] ) );
  DFFX1 \mem_reg[30][28]  ( .D(n1102), .CLK(clk), .Q(\mem[30][28] ) );
  DFFX1 \mem_reg[30][27]  ( .D(n1101), .CLK(clk), .Q(\mem[30][27] ) );
  DFFX1 \mem_reg[30][26]  ( .D(n1100), .CLK(clk), .Q(\mem[30][26] ) );
  DFFX1 \mem_reg[30][25]  ( .D(n1099), .CLK(clk), .Q(\mem[30][25] ) );
  DFFX1 \mem_reg[30][24]  ( .D(n1098), .CLK(clk), .Q(\mem[30][24] ) );
  DFFX1 \mem_reg[30][23]  ( .D(n1097), .CLK(clk), .Q(\mem[30][23] ) );
  DFFX1 \mem_reg[30][22]  ( .D(n1096), .CLK(clk), .Q(\mem[30][22] ) );
  DFFX1 \mem_reg[30][21]  ( .D(n1095), .CLK(clk), .Q(\mem[30][21] ) );
  DFFX1 \mem_reg[30][20]  ( .D(n1094), .CLK(clk), .Q(\mem[30][20] ) );
  DFFX1 \mem_reg[30][19]  ( .D(n1093), .CLK(clk), .Q(\mem[30][19] ) );
  DFFX1 \mem_reg[30][18]  ( .D(n1092), .CLK(clk), .Q(\mem[30][18] ) );
  DFFX1 \mem_reg[30][17]  ( .D(n1091), .CLK(clk), .Q(\mem[30][17] ) );
  DFFX1 \mem_reg[30][16]  ( .D(n1090), .CLK(clk), .Q(\mem[30][16] ) );
  DFFX1 \mem_reg[30][15]  ( .D(n1089), .CLK(clk), .Q(\mem[30][15] ) );
  DFFX1 \mem_reg[30][14]  ( .D(n1088), .CLK(clk), .Q(\mem[30][14] ) );
  DFFX1 \mem_reg[30][13]  ( .D(n1087), .CLK(clk), .Q(\mem[30][13] ) );
  DFFX1 \mem_reg[30][12]  ( .D(n1086), .CLK(clk), .Q(\mem[30][12] ) );
  DFFX1 \mem_reg[30][11]  ( .D(n1085), .CLK(clk), .Q(\mem[30][11] ) );
  DFFX1 \mem_reg[30][10]  ( .D(n1084), .CLK(clk), .Q(\mem[30][10] ) );
  DFFX1 \mem_reg[30][9]  ( .D(n1083), .CLK(clk), .Q(\mem[30][9] ) );
  DFFX1 \mem_reg[30][8]  ( .D(n1082), .CLK(clk), .Q(\mem[30][8] ) );
  DFFX1 \mem_reg[30][7]  ( .D(n1081), .CLK(clk), .Q(\mem[30][7] ) );
  DFFX1 \mem_reg[30][6]  ( .D(n1080), .CLK(clk), .Q(\mem[30][6] ) );
  DFFX1 \mem_reg[30][5]  ( .D(n1079), .CLK(clk), .Q(\mem[30][5] ) );
  DFFX1 \mem_reg[30][4]  ( .D(n1078), .CLK(clk), .Q(\mem[30][4] ) );
  DFFX1 \mem_reg[30][3]  ( .D(n1077), .CLK(clk), .Q(\mem[30][3] ) );
  DFFX1 \mem_reg[30][2]  ( .D(n1076), .CLK(clk), .Q(\mem[30][2] ) );
  DFFX1 \mem_reg[30][1]  ( .D(n1075), .CLK(clk), .Q(\mem[30][1] ) );
  DFFX1 \mem_reg[30][0]  ( .D(n1074), .CLK(clk), .Q(\mem[30][0] ) );
  DFFX1 \mem_reg[29][31]  ( .D(n1073), .CLK(clk), .Q(\mem[29][31] ) );
  DFFX1 \mem_reg[29][30]  ( .D(n1072), .CLK(clk), .Q(\mem[29][30] ) );
  DFFX1 \mem_reg[29][29]  ( .D(n1071), .CLK(clk), .Q(\mem[29][29] ) );
  DFFX1 \mem_reg[29][28]  ( .D(n1070), .CLK(clk), .Q(\mem[29][28] ) );
  DFFX1 \mem_reg[29][27]  ( .D(n1069), .CLK(clk), .Q(\mem[29][27] ) );
  DFFX1 \mem_reg[29][26]  ( .D(n1068), .CLK(clk), .Q(\mem[29][26] ) );
  DFFX1 \mem_reg[29][25]  ( .D(n1067), .CLK(clk), .Q(\mem[29][25] ) );
  DFFX1 \mem_reg[29][24]  ( .D(n1066), .CLK(clk), .Q(\mem[29][24] ) );
  DFFX1 \mem_reg[29][23]  ( .D(n1065), .CLK(clk), .Q(\mem[29][23] ) );
  DFFX1 \mem_reg[29][22]  ( .D(n1064), .CLK(clk), .Q(\mem[29][22] ) );
  DFFX1 \mem_reg[29][21]  ( .D(n1063), .CLK(clk), .Q(\mem[29][21] ) );
  DFFX1 \mem_reg[29][20]  ( .D(n1062), .CLK(clk), .Q(\mem[29][20] ) );
  DFFX1 \mem_reg[29][19]  ( .D(n1061), .CLK(clk), .Q(\mem[29][19] ) );
  DFFX1 \mem_reg[29][18]  ( .D(n1060), .CLK(clk), .Q(\mem[29][18] ) );
  DFFX1 \mem_reg[29][17]  ( .D(n1059), .CLK(clk), .Q(\mem[29][17] ) );
  DFFX1 \mem_reg[29][16]  ( .D(n1058), .CLK(clk), .Q(\mem[29][16] ) );
  DFFX1 \mem_reg[29][15]  ( .D(n1057), .CLK(clk), .Q(\mem[29][15] ) );
  DFFX1 \mem_reg[29][14]  ( .D(n1056), .CLK(clk), .Q(\mem[29][14] ) );
  DFFX1 \mem_reg[29][13]  ( .D(n1055), .CLK(clk), .Q(\mem[29][13] ) );
  DFFX1 \mem_reg[29][12]  ( .D(n1054), .CLK(clk), .Q(\mem[29][12] ) );
  DFFX1 \mem_reg[29][11]  ( .D(n1053), .CLK(clk), .Q(\mem[29][11] ) );
  DFFX1 \mem_reg[29][10]  ( .D(n1052), .CLK(clk), .Q(\mem[29][10] ) );
  DFFX1 \mem_reg[29][9]  ( .D(n1051), .CLK(clk), .Q(\mem[29][9] ) );
  DFFX1 \mem_reg[29][8]  ( .D(n1050), .CLK(clk), .Q(\mem[29][8] ) );
  DFFX1 \mem_reg[29][7]  ( .D(n1049), .CLK(clk), .Q(\mem[29][7] ) );
  DFFX1 \mem_reg[29][6]  ( .D(n1048), .CLK(clk), .Q(\mem[29][6] ) );
  DFFX1 \mem_reg[29][5]  ( .D(n1047), .CLK(clk), .Q(\mem[29][5] ) );
  DFFX1 \mem_reg[29][4]  ( .D(n1046), .CLK(clk), .Q(\mem[29][4] ) );
  DFFX1 \mem_reg[29][3]  ( .D(n1045), .CLK(clk), .Q(\mem[29][3] ) );
  DFFX1 \mem_reg[29][2]  ( .D(n1044), .CLK(clk), .Q(\mem[29][2] ) );
  DFFX1 \mem_reg[29][1]  ( .D(n1043), .CLK(clk), .Q(\mem[29][1] ) );
  DFFX1 \mem_reg[29][0]  ( .D(n1042), .CLK(clk), .Q(\mem[29][0] ) );
  DFFX1 \mem_reg[28][31]  ( .D(n1041), .CLK(clk), .Q(\mem[28][31] ) );
  DFFX1 \mem_reg[28][30]  ( .D(n1040), .CLK(clk), .Q(\mem[28][30] ) );
  DFFX1 \mem_reg[28][29]  ( .D(n1039), .CLK(clk), .Q(\mem[28][29] ) );
  DFFX1 \mem_reg[28][28]  ( .D(n1038), .CLK(clk), .Q(\mem[28][28] ) );
  DFFX1 \mem_reg[28][27]  ( .D(n1037), .CLK(clk), .Q(\mem[28][27] ) );
  DFFX1 \mem_reg[28][26]  ( .D(n1036), .CLK(clk), .Q(\mem[28][26] ) );
  DFFX1 \mem_reg[28][25]  ( .D(n1035), .CLK(clk), .Q(\mem[28][25] ) );
  DFFX1 \mem_reg[28][24]  ( .D(n1034), .CLK(clk), .Q(\mem[28][24] ) );
  DFFX1 \mem_reg[28][23]  ( .D(n1033), .CLK(clk), .Q(\mem[28][23] ) );
  DFFX1 \mem_reg[28][22]  ( .D(n1032), .CLK(clk), .Q(\mem[28][22] ) );
  DFFX1 \mem_reg[28][21]  ( .D(n1031), .CLK(clk), .Q(\mem[28][21] ) );
  DFFX1 \mem_reg[28][20]  ( .D(n1030), .CLK(clk), .Q(\mem[28][20] ) );
  DFFX1 \mem_reg[28][19]  ( .D(n1029), .CLK(clk), .Q(\mem[28][19] ) );
  DFFX1 \mem_reg[28][18]  ( .D(n1028), .CLK(clk), .Q(\mem[28][18] ) );
  DFFX1 \mem_reg[28][17]  ( .D(n1027), .CLK(clk), .Q(\mem[28][17] ) );
  DFFX1 \mem_reg[28][16]  ( .D(n1026), .CLK(clk), .Q(\mem[28][16] ) );
  DFFX1 \mem_reg[28][15]  ( .D(n1025), .CLK(clk), .Q(\mem[28][15] ) );
  DFFX1 \mem_reg[28][14]  ( .D(n1024), .CLK(clk), .Q(\mem[28][14] ) );
  DFFX1 \mem_reg[28][13]  ( .D(n1023), .CLK(clk), .Q(\mem[28][13] ) );
  DFFX1 \mem_reg[28][12]  ( .D(n1022), .CLK(clk), .Q(\mem[28][12] ) );
  DFFX1 \mem_reg[28][11]  ( .D(n1021), .CLK(clk), .Q(\mem[28][11] ) );
  DFFX1 \mem_reg[28][10]  ( .D(n1020), .CLK(clk), .Q(\mem[28][10] ) );
  DFFX1 \mem_reg[28][9]  ( .D(n1019), .CLK(clk), .Q(\mem[28][9] ) );
  DFFX1 \mem_reg[28][8]  ( .D(n1018), .CLK(clk), .Q(\mem[28][8] ) );
  DFFX1 \mem_reg[28][7]  ( .D(n1017), .CLK(clk), .Q(\mem[28][7] ) );
  DFFX1 \mem_reg[28][6]  ( .D(n1016), .CLK(clk), .Q(\mem[28][6] ) );
  DFFX1 \mem_reg[28][5]  ( .D(n1015), .CLK(clk), .Q(\mem[28][5] ) );
  DFFX1 \mem_reg[28][4]  ( .D(n1014), .CLK(clk), .Q(\mem[28][4] ) );
  DFFX1 \mem_reg[28][3]  ( .D(n1013), .CLK(clk), .Q(\mem[28][3] ) );
  DFFX1 \mem_reg[28][2]  ( .D(n1012), .CLK(clk), .Q(\mem[28][2] ) );
  DFFX1 \mem_reg[28][1]  ( .D(n1011), .CLK(clk), .Q(\mem[28][1] ) );
  DFFX1 \mem_reg[28][0]  ( .D(n1010), .CLK(clk), .Q(\mem[28][0] ) );
  DFFX1 \mem_reg[27][31]  ( .D(n1009), .CLK(clk), .Q(\mem[27][31] ) );
  DFFX1 \mem_reg[27][30]  ( .D(n1008), .CLK(clk), .Q(\mem[27][30] ) );
  DFFX1 \mem_reg[27][29]  ( .D(n1007), .CLK(clk), .Q(\mem[27][29] ) );
  DFFX1 \mem_reg[27][28]  ( .D(n1006), .CLK(clk), .Q(\mem[27][28] ) );
  DFFX1 \mem_reg[27][27]  ( .D(n1005), .CLK(clk), .Q(\mem[27][27] ) );
  DFFX1 \mem_reg[27][26]  ( .D(n1004), .CLK(clk), .Q(\mem[27][26] ) );
  DFFX1 \mem_reg[27][25]  ( .D(n1003), .CLK(clk), .Q(\mem[27][25] ) );
  DFFX1 \mem_reg[27][24]  ( .D(n1002), .CLK(clk), .Q(\mem[27][24] ) );
  DFFX1 \mem_reg[27][23]  ( .D(n1001), .CLK(clk), .Q(\mem[27][23] ) );
  DFFX1 \mem_reg[27][22]  ( .D(n1000), .CLK(clk), .Q(\mem[27][22] ) );
  DFFX1 \mem_reg[27][21]  ( .D(n999), .CLK(clk), .Q(\mem[27][21] ) );
  DFFX1 \mem_reg[27][20]  ( .D(n998), .CLK(clk), .Q(\mem[27][20] ) );
  DFFX1 \mem_reg[27][19]  ( .D(n997), .CLK(clk), .Q(\mem[27][19] ) );
  DFFX1 \mem_reg[27][18]  ( .D(n996), .CLK(clk), .Q(\mem[27][18] ) );
  DFFX1 \mem_reg[27][17]  ( .D(n995), .CLK(clk), .Q(\mem[27][17] ) );
  DFFX1 \mem_reg[27][16]  ( .D(n994), .CLK(clk), .Q(\mem[27][16] ) );
  DFFX1 \mem_reg[27][15]  ( .D(n993), .CLK(clk), .Q(\mem[27][15] ) );
  DFFX1 \mem_reg[27][14]  ( .D(n992), .CLK(clk), .Q(\mem[27][14] ) );
  DFFX1 \mem_reg[27][13]  ( .D(n991), .CLK(clk), .Q(\mem[27][13] ) );
  DFFX1 \mem_reg[27][12]  ( .D(n990), .CLK(clk), .Q(\mem[27][12] ) );
  DFFX1 \mem_reg[27][11]  ( .D(n989), .CLK(clk), .Q(\mem[27][11] ) );
  DFFX1 \mem_reg[27][10]  ( .D(n988), .CLK(clk), .Q(\mem[27][10] ) );
  DFFX1 \mem_reg[27][9]  ( .D(n987), .CLK(clk), .Q(\mem[27][9] ) );
  DFFX1 \mem_reg[27][8]  ( .D(n986), .CLK(clk), .Q(\mem[27][8] ) );
  DFFX1 \mem_reg[27][7]  ( .D(n985), .CLK(clk), .Q(\mem[27][7] ) );
  DFFX1 \mem_reg[27][6]  ( .D(n984), .CLK(clk), .Q(\mem[27][6] ) );
  DFFX1 \mem_reg[27][5]  ( .D(n983), .CLK(clk), .Q(\mem[27][5] ) );
  DFFX1 \mem_reg[27][4]  ( .D(n982), .CLK(clk), .Q(\mem[27][4] ) );
  DFFX1 \mem_reg[27][3]  ( .D(n981), .CLK(clk), .Q(\mem[27][3] ) );
  DFFX1 \mem_reg[27][2]  ( .D(n980), .CLK(clk), .Q(\mem[27][2] ) );
  DFFX1 \mem_reg[27][1]  ( .D(n979), .CLK(clk), .Q(\mem[27][1] ) );
  DFFX1 \mem_reg[27][0]  ( .D(n978), .CLK(clk), .Q(\mem[27][0] ) );
  DFFX1 \mem_reg[26][31]  ( .D(n977), .CLK(clk), .Q(\mem[26][31] ) );
  DFFX1 \mem_reg[26][30]  ( .D(n976), .CLK(clk), .Q(\mem[26][30] ) );
  DFFX1 \mem_reg[26][29]  ( .D(n975), .CLK(clk), .Q(\mem[26][29] ) );
  DFFX1 \mem_reg[26][28]  ( .D(n974), .CLK(clk), .Q(\mem[26][28] ) );
  DFFX1 \mem_reg[26][27]  ( .D(n973), .CLK(clk), .Q(\mem[26][27] ) );
  DFFX1 \mem_reg[26][26]  ( .D(n972), .CLK(clk), .Q(\mem[26][26] ) );
  DFFX1 \mem_reg[26][25]  ( .D(n971), .CLK(clk), .Q(\mem[26][25] ) );
  DFFX1 \mem_reg[26][24]  ( .D(n970), .CLK(clk), .Q(\mem[26][24] ) );
  DFFX1 \mem_reg[26][23]  ( .D(n969), .CLK(clk), .Q(\mem[26][23] ) );
  DFFX1 \mem_reg[26][22]  ( .D(n968), .CLK(clk), .Q(\mem[26][22] ) );
  DFFX1 \mem_reg[26][21]  ( .D(n967), .CLK(clk), .Q(\mem[26][21] ) );
  DFFX1 \mem_reg[26][20]  ( .D(n966), .CLK(clk), .Q(\mem[26][20] ) );
  DFFX1 \mem_reg[26][19]  ( .D(n965), .CLK(clk), .Q(\mem[26][19] ) );
  DFFX1 \mem_reg[26][18]  ( .D(n964), .CLK(clk), .Q(\mem[26][18] ) );
  DFFX1 \mem_reg[26][17]  ( .D(n963), .CLK(clk), .Q(\mem[26][17] ) );
  DFFX1 \mem_reg[26][16]  ( .D(n962), .CLK(clk), .Q(\mem[26][16] ) );
  DFFX1 \mem_reg[26][15]  ( .D(n961), .CLK(clk), .Q(\mem[26][15] ) );
  DFFX1 \mem_reg[26][14]  ( .D(n960), .CLK(clk), .Q(\mem[26][14] ) );
  DFFX1 \mem_reg[26][13]  ( .D(n959), .CLK(clk), .Q(\mem[26][13] ) );
  DFFX1 \mem_reg[26][12]  ( .D(n958), .CLK(clk), .Q(\mem[26][12] ) );
  DFFX1 \mem_reg[26][11]  ( .D(n957), .CLK(clk), .Q(\mem[26][11] ) );
  DFFX1 \mem_reg[26][10]  ( .D(n956), .CLK(clk), .Q(\mem[26][10] ) );
  DFFX1 \mem_reg[26][9]  ( .D(n955), .CLK(clk), .Q(\mem[26][9] ) );
  DFFX1 \mem_reg[26][8]  ( .D(n954), .CLK(clk), .Q(\mem[26][8] ) );
  DFFX1 \mem_reg[26][7]  ( .D(n953), .CLK(clk), .Q(\mem[26][7] ) );
  DFFX1 \mem_reg[26][6]  ( .D(n952), .CLK(clk), .Q(\mem[26][6] ) );
  DFFX1 \mem_reg[26][5]  ( .D(n951), .CLK(clk), .Q(\mem[26][5] ) );
  DFFX1 \mem_reg[26][4]  ( .D(n950), .CLK(clk), .Q(\mem[26][4] ) );
  DFFX1 \mem_reg[26][3]  ( .D(n949), .CLK(clk), .Q(\mem[26][3] ) );
  DFFX1 \mem_reg[26][2]  ( .D(n948), .CLK(clk), .Q(\mem[26][2] ) );
  DFFX1 \mem_reg[26][1]  ( .D(n947), .CLK(clk), .Q(\mem[26][1] ) );
  DFFX1 \mem_reg[26][0]  ( .D(n946), .CLK(clk), .Q(\mem[26][0] ) );
  DFFX1 \mem_reg[25][31]  ( .D(n945), .CLK(clk), .Q(\mem[25][31] ) );
  DFFX1 \mem_reg[25][30]  ( .D(n944), .CLK(clk), .Q(\mem[25][30] ) );
  DFFX1 \mem_reg[25][29]  ( .D(n943), .CLK(clk), .Q(\mem[25][29] ) );
  DFFX1 \mem_reg[25][28]  ( .D(n942), .CLK(clk), .Q(\mem[25][28] ) );
  DFFX1 \mem_reg[25][27]  ( .D(n941), .CLK(clk), .Q(\mem[25][27] ) );
  DFFX1 \mem_reg[25][26]  ( .D(n940), .CLK(clk), .Q(\mem[25][26] ) );
  DFFX1 \mem_reg[25][25]  ( .D(n939), .CLK(clk), .Q(\mem[25][25] ) );
  DFFX1 \mem_reg[25][24]  ( .D(n938), .CLK(clk), .Q(\mem[25][24] ) );
  DFFX1 \mem_reg[25][23]  ( .D(n937), .CLK(clk), .Q(\mem[25][23] ) );
  DFFX1 \mem_reg[25][22]  ( .D(n936), .CLK(clk), .Q(\mem[25][22] ) );
  DFFX1 \mem_reg[25][21]  ( .D(n935), .CLK(clk), .Q(\mem[25][21] ) );
  DFFX1 \mem_reg[25][20]  ( .D(n934), .CLK(clk), .Q(\mem[25][20] ) );
  DFFX1 \mem_reg[25][19]  ( .D(n933), .CLK(clk), .Q(\mem[25][19] ) );
  DFFX1 \mem_reg[25][18]  ( .D(n932), .CLK(clk), .Q(\mem[25][18] ) );
  DFFX1 \mem_reg[25][17]  ( .D(n931), .CLK(clk), .Q(\mem[25][17] ) );
  DFFX1 \mem_reg[25][16]  ( .D(n930), .CLK(clk), .Q(\mem[25][16] ) );
  DFFX1 \mem_reg[25][15]  ( .D(n929), .CLK(clk), .Q(\mem[25][15] ) );
  DFFX1 \mem_reg[25][14]  ( .D(n928), .CLK(clk), .Q(\mem[25][14] ) );
  DFFX1 \mem_reg[25][13]  ( .D(n927), .CLK(clk), .Q(\mem[25][13] ) );
  DFFX1 \mem_reg[25][12]  ( .D(n926), .CLK(clk), .Q(\mem[25][12] ) );
  DFFX1 \mem_reg[25][11]  ( .D(n925), .CLK(clk), .Q(\mem[25][11] ) );
  DFFX1 \mem_reg[25][10]  ( .D(n924), .CLK(clk), .Q(\mem[25][10] ) );
  DFFX1 \mem_reg[25][9]  ( .D(n923), .CLK(clk), .Q(\mem[25][9] ) );
  DFFX1 \mem_reg[25][8]  ( .D(n922), .CLK(clk), .Q(\mem[25][8] ) );
  DFFX1 \mem_reg[25][7]  ( .D(n921), .CLK(clk), .Q(\mem[25][7] ) );
  DFFX1 \mem_reg[25][6]  ( .D(n920), .CLK(clk), .Q(\mem[25][6] ) );
  DFFX1 \mem_reg[25][5]  ( .D(n919), .CLK(clk), .Q(\mem[25][5] ) );
  DFFX1 \mem_reg[25][4]  ( .D(n918), .CLK(clk), .Q(\mem[25][4] ) );
  DFFX1 \mem_reg[25][3]  ( .D(n917), .CLK(clk), .Q(\mem[25][3] ) );
  DFFX1 \mem_reg[25][2]  ( .D(n916), .CLK(clk), .Q(\mem[25][2] ) );
  DFFX1 \mem_reg[25][1]  ( .D(n915), .CLK(clk), .Q(\mem[25][1] ) );
  DFFX1 \mem_reg[25][0]  ( .D(n914), .CLK(clk), .Q(\mem[25][0] ) );
  DFFX1 \mem_reg[24][31]  ( .D(n913), .CLK(clk), .Q(\mem[24][31] ) );
  DFFX1 \mem_reg[24][30]  ( .D(n912), .CLK(clk), .Q(\mem[24][30] ) );
  DFFX1 \mem_reg[24][29]  ( .D(n911), .CLK(clk), .Q(\mem[24][29] ) );
  DFFX1 \mem_reg[24][28]  ( .D(n910), .CLK(clk), .Q(\mem[24][28] ) );
  DFFX1 \mem_reg[24][27]  ( .D(n909), .CLK(clk), .Q(\mem[24][27] ) );
  DFFX1 \mem_reg[24][26]  ( .D(n908), .CLK(clk), .Q(\mem[24][26] ) );
  DFFX1 \mem_reg[24][25]  ( .D(n907), .CLK(clk), .Q(\mem[24][25] ) );
  DFFX1 \mem_reg[24][24]  ( .D(n906), .CLK(clk), .Q(\mem[24][24] ) );
  DFFX1 \mem_reg[24][23]  ( .D(n905), .CLK(clk), .Q(\mem[24][23] ) );
  DFFX1 \mem_reg[24][22]  ( .D(n904), .CLK(clk), .Q(\mem[24][22] ) );
  DFFX1 \mem_reg[24][21]  ( .D(n903), .CLK(clk), .Q(\mem[24][21] ) );
  DFFX1 \mem_reg[24][20]  ( .D(n902), .CLK(clk), .Q(\mem[24][20] ) );
  DFFX1 \mem_reg[24][19]  ( .D(n901), .CLK(clk), .Q(\mem[24][19] ) );
  DFFX1 \mem_reg[24][18]  ( .D(n900), .CLK(clk), .Q(\mem[24][18] ) );
  DFFX1 \mem_reg[24][17]  ( .D(n899), .CLK(clk), .Q(\mem[24][17] ) );
  DFFX1 \mem_reg[24][16]  ( .D(n898), .CLK(clk), .Q(\mem[24][16] ) );
  DFFX1 \mem_reg[24][15]  ( .D(n897), .CLK(clk), .Q(\mem[24][15] ) );
  DFFX1 \mem_reg[24][14]  ( .D(n896), .CLK(clk), .Q(\mem[24][14] ) );
  DFFX1 \mem_reg[24][13]  ( .D(n895), .CLK(clk), .Q(\mem[24][13] ) );
  DFFX1 \mem_reg[24][12]  ( .D(n894), .CLK(clk), .Q(\mem[24][12] ) );
  DFFX1 \mem_reg[24][11]  ( .D(n893), .CLK(clk), .Q(\mem[24][11] ) );
  DFFX1 \mem_reg[24][10]  ( .D(n892), .CLK(clk), .Q(\mem[24][10] ) );
  DFFX1 \mem_reg[24][9]  ( .D(n891), .CLK(clk), .Q(\mem[24][9] ) );
  DFFX1 \mem_reg[24][8]  ( .D(n890), .CLK(clk), .Q(\mem[24][8] ) );
  DFFX1 \mem_reg[24][7]  ( .D(n889), .CLK(clk), .Q(\mem[24][7] ) );
  DFFX1 \mem_reg[24][6]  ( .D(n888), .CLK(clk), .Q(\mem[24][6] ) );
  DFFX1 \mem_reg[24][5]  ( .D(n887), .CLK(clk), .Q(\mem[24][5] ) );
  DFFX1 \mem_reg[24][4]  ( .D(n886), .CLK(clk), .Q(\mem[24][4] ) );
  DFFX1 \mem_reg[24][3]  ( .D(n885), .CLK(clk), .Q(\mem[24][3] ) );
  DFFX1 \mem_reg[24][2]  ( .D(n884), .CLK(clk), .Q(\mem[24][2] ) );
  DFFX1 \mem_reg[24][1]  ( .D(n883), .CLK(clk), .Q(\mem[24][1] ) );
  DFFX1 \mem_reg[24][0]  ( .D(n882), .CLK(clk), .Q(\mem[24][0] ) );
  DFFX1 \mem_reg[23][31]  ( .D(n881), .CLK(clk), .Q(\mem[23][31] ) );
  DFFX1 \mem_reg[23][30]  ( .D(n880), .CLK(clk), .Q(\mem[23][30] ) );
  DFFX1 \mem_reg[23][29]  ( .D(n879), .CLK(clk), .Q(\mem[23][29] ) );
  DFFX1 \mem_reg[23][28]  ( .D(n878), .CLK(clk), .Q(\mem[23][28] ) );
  DFFX1 \mem_reg[23][27]  ( .D(n877), .CLK(clk), .Q(\mem[23][27] ) );
  DFFX1 \mem_reg[23][26]  ( .D(n876), .CLK(clk), .Q(\mem[23][26] ) );
  DFFX1 \mem_reg[23][25]  ( .D(n875), .CLK(clk), .Q(\mem[23][25] ) );
  DFFX1 \mem_reg[23][24]  ( .D(n874), .CLK(clk), .Q(\mem[23][24] ) );
  DFFX1 \mem_reg[23][23]  ( .D(n873), .CLK(clk), .Q(\mem[23][23] ) );
  DFFX1 \mem_reg[23][22]  ( .D(n872), .CLK(clk), .Q(\mem[23][22] ) );
  DFFX1 \mem_reg[23][21]  ( .D(n871), .CLK(clk), .Q(\mem[23][21] ) );
  DFFX1 \mem_reg[23][20]  ( .D(n870), .CLK(clk), .Q(\mem[23][20] ) );
  DFFX1 \mem_reg[23][19]  ( .D(n869), .CLK(clk), .Q(\mem[23][19] ) );
  DFFX1 \mem_reg[23][18]  ( .D(n868), .CLK(clk), .Q(\mem[23][18] ) );
  DFFX1 \mem_reg[23][17]  ( .D(n867), .CLK(clk), .Q(\mem[23][17] ) );
  DFFX1 \mem_reg[23][16]  ( .D(n866), .CLK(clk), .Q(\mem[23][16] ) );
  DFFX1 \mem_reg[23][15]  ( .D(n865), .CLK(clk), .Q(\mem[23][15] ) );
  DFFX1 \mem_reg[23][14]  ( .D(n864), .CLK(clk), .Q(\mem[23][14] ) );
  DFFX1 \mem_reg[23][13]  ( .D(n863), .CLK(clk), .Q(\mem[23][13] ) );
  DFFX1 \mem_reg[23][12]  ( .D(n862), .CLK(clk), .Q(\mem[23][12] ) );
  DFFX1 \mem_reg[23][11]  ( .D(n861), .CLK(clk), .Q(\mem[23][11] ) );
  DFFX1 \mem_reg[23][10]  ( .D(n860), .CLK(clk), .Q(\mem[23][10] ) );
  DFFX1 \mem_reg[23][9]  ( .D(n859), .CLK(clk), .Q(\mem[23][9] ) );
  DFFX1 \mem_reg[23][8]  ( .D(n858), .CLK(clk), .Q(\mem[23][8] ) );
  DFFX1 \mem_reg[23][7]  ( .D(n857), .CLK(clk), .Q(\mem[23][7] ) );
  DFFX1 \mem_reg[23][6]  ( .D(n856), .CLK(clk), .Q(\mem[23][6] ) );
  DFFX1 \mem_reg[23][5]  ( .D(n855), .CLK(clk), .Q(\mem[23][5] ) );
  DFFX1 \mem_reg[23][4]  ( .D(n854), .CLK(clk), .Q(\mem[23][4] ) );
  DFFX1 \mem_reg[23][3]  ( .D(n853), .CLK(clk), .Q(\mem[23][3] ) );
  DFFX1 \mem_reg[23][2]  ( .D(n852), .CLK(clk), .Q(\mem[23][2] ) );
  DFFX1 \mem_reg[23][1]  ( .D(n851), .CLK(clk), .Q(\mem[23][1] ) );
  DFFX1 \mem_reg[23][0]  ( .D(n850), .CLK(clk), .Q(\mem[23][0] ) );
  DFFX1 \mem_reg[22][31]  ( .D(n849), .CLK(clk), .Q(\mem[22][31] ) );
  DFFX1 \mem_reg[22][30]  ( .D(n848), .CLK(clk), .Q(\mem[22][30] ) );
  DFFX1 \mem_reg[22][29]  ( .D(n847), .CLK(clk), .Q(\mem[22][29] ) );
  DFFX1 \mem_reg[22][28]  ( .D(n846), .CLK(clk), .Q(\mem[22][28] ) );
  DFFX1 \mem_reg[22][27]  ( .D(n845), .CLK(clk), .Q(\mem[22][27] ) );
  DFFX1 \mem_reg[22][26]  ( .D(n844), .CLK(clk), .Q(\mem[22][26] ) );
  DFFX1 \mem_reg[22][25]  ( .D(n843), .CLK(clk), .Q(\mem[22][25] ) );
  DFFX1 \mem_reg[22][24]  ( .D(n842), .CLK(clk), .Q(\mem[22][24] ) );
  DFFX1 \mem_reg[22][23]  ( .D(n841), .CLK(clk), .Q(\mem[22][23] ) );
  DFFX1 \mem_reg[22][22]  ( .D(n840), .CLK(clk), .Q(\mem[22][22] ) );
  DFFX1 \mem_reg[22][21]  ( .D(n839), .CLK(clk), .Q(\mem[22][21] ) );
  DFFX1 \mem_reg[22][20]  ( .D(n838), .CLK(clk), .Q(\mem[22][20] ) );
  DFFX1 \mem_reg[22][19]  ( .D(n837), .CLK(clk), .Q(\mem[22][19] ) );
  DFFX1 \mem_reg[22][18]  ( .D(n836), .CLK(clk), .Q(\mem[22][18] ) );
  DFFX1 \mem_reg[22][17]  ( .D(n835), .CLK(clk), .Q(\mem[22][17] ) );
  DFFX1 \mem_reg[22][16]  ( .D(n834), .CLK(clk), .Q(\mem[22][16] ) );
  DFFX1 \mem_reg[22][15]  ( .D(n833), .CLK(clk), .Q(\mem[22][15] ) );
  DFFX1 \mem_reg[22][14]  ( .D(n832), .CLK(clk), .Q(\mem[22][14] ) );
  DFFX1 \mem_reg[22][13]  ( .D(n831), .CLK(clk), .Q(\mem[22][13] ) );
  DFFX1 \mem_reg[22][12]  ( .D(n830), .CLK(clk), .Q(\mem[22][12] ) );
  DFFX1 \mem_reg[22][11]  ( .D(n829), .CLK(clk), .Q(\mem[22][11] ) );
  DFFX1 \mem_reg[22][10]  ( .D(n828), .CLK(clk), .Q(\mem[22][10] ) );
  DFFX1 \mem_reg[22][9]  ( .D(n827), .CLK(clk), .Q(\mem[22][9] ) );
  DFFX1 \mem_reg[22][8]  ( .D(n826), .CLK(clk), .Q(\mem[22][8] ) );
  DFFX1 \mem_reg[22][7]  ( .D(n825), .CLK(clk), .Q(\mem[22][7] ) );
  DFFX1 \mem_reg[22][6]  ( .D(n824), .CLK(clk), .Q(\mem[22][6] ) );
  DFFX1 \mem_reg[22][5]  ( .D(n823), .CLK(clk), .Q(\mem[22][5] ) );
  DFFX1 \mem_reg[22][4]  ( .D(n822), .CLK(clk), .Q(\mem[22][4] ) );
  DFFX1 \mem_reg[22][3]  ( .D(n821), .CLK(clk), .Q(\mem[22][3] ) );
  DFFX1 \mem_reg[22][2]  ( .D(n820), .CLK(clk), .Q(\mem[22][2] ) );
  DFFX1 \mem_reg[22][1]  ( .D(n819), .CLK(clk), .Q(\mem[22][1] ) );
  DFFX1 \mem_reg[22][0]  ( .D(n818), .CLK(clk), .Q(\mem[22][0] ) );
  DFFX1 \mem_reg[21][31]  ( .D(n817), .CLK(clk), .Q(\mem[21][31] ) );
  DFFX1 \mem_reg[21][30]  ( .D(n816), .CLK(clk), .Q(\mem[21][30] ) );
  DFFX1 \mem_reg[21][29]  ( .D(n815), .CLK(clk), .Q(\mem[21][29] ) );
  DFFX1 \mem_reg[21][28]  ( .D(n814), .CLK(clk), .Q(\mem[21][28] ) );
  DFFX1 \mem_reg[21][27]  ( .D(n813), .CLK(clk), .Q(\mem[21][27] ) );
  DFFX1 \mem_reg[21][26]  ( .D(n812), .CLK(clk), .Q(\mem[21][26] ) );
  DFFX1 \mem_reg[21][25]  ( .D(n811), .CLK(clk), .Q(\mem[21][25] ) );
  DFFX1 \mem_reg[21][24]  ( .D(n810), .CLK(clk), .Q(\mem[21][24] ) );
  DFFX1 \mem_reg[21][23]  ( .D(n809), .CLK(clk), .Q(\mem[21][23] ) );
  DFFX1 \mem_reg[21][22]  ( .D(n808), .CLK(clk), .Q(\mem[21][22] ) );
  DFFX1 \mem_reg[21][21]  ( .D(n807), .CLK(clk), .Q(\mem[21][21] ) );
  DFFX1 \mem_reg[21][20]  ( .D(n806), .CLK(clk), .Q(\mem[21][20] ) );
  DFFX1 \mem_reg[21][19]  ( .D(n805), .CLK(clk), .Q(\mem[21][19] ) );
  DFFX1 \mem_reg[21][18]  ( .D(n804), .CLK(clk), .Q(\mem[21][18] ) );
  DFFX1 \mem_reg[21][17]  ( .D(n803), .CLK(clk), .Q(\mem[21][17] ) );
  DFFX1 \mem_reg[21][16]  ( .D(n802), .CLK(clk), .Q(\mem[21][16] ) );
  DFFX1 \mem_reg[21][15]  ( .D(n801), .CLK(clk), .Q(\mem[21][15] ) );
  DFFX1 \mem_reg[21][14]  ( .D(n800), .CLK(clk), .Q(\mem[21][14] ) );
  DFFX1 \mem_reg[21][13]  ( .D(n799), .CLK(clk), .Q(\mem[21][13] ) );
  DFFX1 \mem_reg[21][12]  ( .D(n798), .CLK(clk), .Q(\mem[21][12] ) );
  DFFX1 \mem_reg[21][11]  ( .D(n797), .CLK(clk), .Q(\mem[21][11] ) );
  DFFX1 \mem_reg[21][10]  ( .D(n796), .CLK(clk), .Q(\mem[21][10] ) );
  DFFX1 \mem_reg[21][9]  ( .D(n795), .CLK(clk), .Q(\mem[21][9] ) );
  DFFX1 \mem_reg[21][8]  ( .D(n794), .CLK(clk), .Q(\mem[21][8] ) );
  DFFX1 \mem_reg[21][7]  ( .D(n793), .CLK(clk), .Q(\mem[21][7] ) );
  DFFX1 \mem_reg[21][6]  ( .D(n792), .CLK(clk), .Q(\mem[21][6] ) );
  DFFX1 \mem_reg[21][5]  ( .D(n791), .CLK(clk), .Q(\mem[21][5] ) );
  DFFX1 \mem_reg[21][4]  ( .D(n790), .CLK(clk), .Q(\mem[21][4] ) );
  DFFX1 \mem_reg[21][3]  ( .D(n789), .CLK(clk), .Q(\mem[21][3] ) );
  DFFX1 \mem_reg[21][2]  ( .D(n788), .CLK(clk), .Q(\mem[21][2] ) );
  DFFX1 \mem_reg[21][1]  ( .D(n787), .CLK(clk), .Q(\mem[21][1] ) );
  DFFX1 \mem_reg[21][0]  ( .D(n786), .CLK(clk), .Q(\mem[21][0] ) );
  DFFX1 \mem_reg[20][31]  ( .D(n785), .CLK(clk), .Q(\mem[20][31] ) );
  DFFX1 \mem_reg[20][30]  ( .D(n784), .CLK(clk), .Q(\mem[20][30] ) );
  DFFX1 \mem_reg[20][29]  ( .D(n783), .CLK(clk), .Q(\mem[20][29] ) );
  DFFX1 \mem_reg[20][28]  ( .D(n782), .CLK(clk), .Q(\mem[20][28] ) );
  DFFX1 \mem_reg[20][27]  ( .D(n781), .CLK(clk), .Q(\mem[20][27] ) );
  DFFX1 \mem_reg[20][26]  ( .D(n780), .CLK(clk), .Q(\mem[20][26] ) );
  DFFX1 \mem_reg[20][25]  ( .D(n779), .CLK(clk), .Q(\mem[20][25] ) );
  DFFX1 \mem_reg[20][24]  ( .D(n778), .CLK(clk), .Q(\mem[20][24] ) );
  DFFX1 \mem_reg[20][23]  ( .D(n777), .CLK(clk), .Q(\mem[20][23] ) );
  DFFX1 \mem_reg[20][22]  ( .D(n776), .CLK(clk), .Q(\mem[20][22] ) );
  DFFX1 \mem_reg[20][21]  ( .D(n775), .CLK(clk), .Q(\mem[20][21] ) );
  DFFX1 \mem_reg[20][20]  ( .D(n774), .CLK(clk), .Q(\mem[20][20] ) );
  DFFX1 \mem_reg[20][19]  ( .D(n773), .CLK(clk), .Q(\mem[20][19] ) );
  DFFX1 \mem_reg[20][18]  ( .D(n772), .CLK(clk), .Q(\mem[20][18] ) );
  DFFX1 \mem_reg[20][17]  ( .D(n771), .CLK(clk), .Q(\mem[20][17] ) );
  DFFX1 \mem_reg[20][16]  ( .D(n770), .CLK(clk), .Q(\mem[20][16] ) );
  DFFX1 \mem_reg[20][15]  ( .D(n769), .CLK(clk), .Q(\mem[20][15] ) );
  DFFX1 \mem_reg[20][14]  ( .D(n768), .CLK(clk), .Q(\mem[20][14] ) );
  DFFX1 \mem_reg[20][13]  ( .D(n767), .CLK(clk), .Q(\mem[20][13] ) );
  DFFX1 \mem_reg[20][12]  ( .D(n766), .CLK(clk), .Q(\mem[20][12] ) );
  DFFX1 \mem_reg[20][11]  ( .D(n765), .CLK(clk), .Q(\mem[20][11] ) );
  DFFX1 \mem_reg[20][10]  ( .D(n764), .CLK(clk), .Q(\mem[20][10] ) );
  DFFX1 \mem_reg[20][9]  ( .D(n763), .CLK(clk), .Q(\mem[20][9] ) );
  DFFX1 \mem_reg[20][8]  ( .D(n762), .CLK(clk), .Q(\mem[20][8] ) );
  DFFX1 \mem_reg[20][7]  ( .D(n761), .CLK(clk), .Q(\mem[20][7] ) );
  DFFX1 \mem_reg[20][6]  ( .D(n760), .CLK(clk), .Q(\mem[20][6] ) );
  DFFX1 \mem_reg[20][5]  ( .D(n759), .CLK(clk), .Q(\mem[20][5] ) );
  DFFX1 \mem_reg[20][4]  ( .D(n758), .CLK(clk), .Q(\mem[20][4] ) );
  DFFX1 \mem_reg[20][3]  ( .D(n757), .CLK(clk), .Q(\mem[20][3] ) );
  DFFX1 \mem_reg[20][2]  ( .D(n756), .CLK(clk), .Q(\mem[20][2] ) );
  DFFX1 \mem_reg[20][1]  ( .D(n755), .CLK(clk), .Q(\mem[20][1] ) );
  DFFX1 \mem_reg[20][0]  ( .D(n754), .CLK(clk), .Q(\mem[20][0] ) );
  DFFX1 \mem_reg[19][31]  ( .D(n753), .CLK(clk), .Q(\mem[19][31] ) );
  DFFX1 \mem_reg[19][30]  ( .D(n752), .CLK(clk), .Q(\mem[19][30] ) );
  DFFX1 \mem_reg[19][29]  ( .D(n751), .CLK(clk), .Q(\mem[19][29] ) );
  DFFX1 \mem_reg[19][28]  ( .D(n750), .CLK(clk), .Q(\mem[19][28] ) );
  DFFX1 \mem_reg[19][27]  ( .D(n749), .CLK(clk), .Q(\mem[19][27] ) );
  DFFX1 \mem_reg[19][26]  ( .D(n748), .CLK(clk), .Q(\mem[19][26] ) );
  DFFX1 \mem_reg[19][25]  ( .D(n747), .CLK(clk), .Q(\mem[19][25] ) );
  DFFX1 \mem_reg[19][24]  ( .D(n746), .CLK(clk), .Q(\mem[19][24] ) );
  DFFX1 \mem_reg[19][23]  ( .D(n745), .CLK(clk), .Q(\mem[19][23] ) );
  DFFX1 \mem_reg[19][22]  ( .D(n744), .CLK(clk), .Q(\mem[19][22] ) );
  DFFX1 \mem_reg[19][21]  ( .D(n743), .CLK(clk), .Q(\mem[19][21] ) );
  DFFX1 \mem_reg[19][20]  ( .D(n742), .CLK(clk), .Q(\mem[19][20] ) );
  DFFX1 \mem_reg[19][19]  ( .D(n741), .CLK(clk), .Q(\mem[19][19] ) );
  DFFX1 \mem_reg[19][18]  ( .D(n740), .CLK(clk), .Q(\mem[19][18] ) );
  DFFX1 \mem_reg[19][17]  ( .D(n739), .CLK(clk), .Q(\mem[19][17] ) );
  DFFX1 \mem_reg[19][16]  ( .D(n738), .CLK(clk), .Q(\mem[19][16] ) );
  DFFX1 \mem_reg[19][15]  ( .D(n737), .CLK(clk), .Q(\mem[19][15] ) );
  DFFX1 \mem_reg[19][14]  ( .D(n736), .CLK(clk), .Q(\mem[19][14] ) );
  DFFX1 \mem_reg[19][13]  ( .D(n735), .CLK(clk), .Q(\mem[19][13] ) );
  DFFX1 \mem_reg[19][12]  ( .D(n734), .CLK(clk), .Q(\mem[19][12] ) );
  DFFX1 \mem_reg[19][11]  ( .D(n733), .CLK(clk), .Q(\mem[19][11] ) );
  DFFX1 \mem_reg[19][10]  ( .D(n732), .CLK(clk), .Q(\mem[19][10] ) );
  DFFX1 \mem_reg[19][9]  ( .D(n731), .CLK(clk), .Q(\mem[19][9] ) );
  DFFX1 \mem_reg[19][8]  ( .D(n730), .CLK(clk), .Q(\mem[19][8] ) );
  DFFX1 \mem_reg[19][7]  ( .D(n729), .CLK(clk), .Q(\mem[19][7] ) );
  DFFX1 \mem_reg[19][6]  ( .D(n728), .CLK(clk), .Q(\mem[19][6] ) );
  DFFX1 \mem_reg[19][5]  ( .D(n727), .CLK(clk), .Q(\mem[19][5] ) );
  DFFX1 \mem_reg[19][4]  ( .D(n726), .CLK(clk), .Q(\mem[19][4] ) );
  DFFX1 \mem_reg[19][3]  ( .D(n725), .CLK(clk), .Q(\mem[19][3] ) );
  DFFX1 \mem_reg[19][2]  ( .D(n724), .CLK(clk), .Q(\mem[19][2] ) );
  DFFX1 \mem_reg[19][1]  ( .D(n723), .CLK(clk), .Q(\mem[19][1] ) );
  DFFX1 \mem_reg[19][0]  ( .D(n722), .CLK(clk), .Q(\mem[19][0] ) );
  DFFX1 \mem_reg[18][31]  ( .D(n721), .CLK(clk), .Q(\mem[18][31] ) );
  DFFX1 \mem_reg[18][30]  ( .D(n720), .CLK(clk), .Q(\mem[18][30] ) );
  DFFX1 \mem_reg[18][29]  ( .D(n719), .CLK(clk), .Q(\mem[18][29] ) );
  DFFX1 \mem_reg[18][28]  ( .D(n718), .CLK(clk), .Q(\mem[18][28] ) );
  DFFX1 \mem_reg[18][27]  ( .D(n717), .CLK(clk), .Q(\mem[18][27] ) );
  DFFX1 \mem_reg[18][26]  ( .D(n716), .CLK(clk), .Q(\mem[18][26] ) );
  DFFX1 \mem_reg[18][25]  ( .D(n715), .CLK(clk), .Q(\mem[18][25] ) );
  DFFX1 \mem_reg[18][24]  ( .D(n714), .CLK(clk), .Q(\mem[18][24] ) );
  DFFX1 \mem_reg[18][23]  ( .D(n713), .CLK(clk), .Q(\mem[18][23] ) );
  DFFX1 \mem_reg[18][22]  ( .D(n712), .CLK(clk), .Q(\mem[18][22] ) );
  DFFX1 \mem_reg[18][21]  ( .D(n711), .CLK(clk), .Q(\mem[18][21] ) );
  DFFX1 \mem_reg[18][20]  ( .D(n710), .CLK(clk), .Q(\mem[18][20] ) );
  DFFX1 \mem_reg[18][19]  ( .D(n709), .CLK(clk), .Q(\mem[18][19] ) );
  DFFX1 \mem_reg[18][18]  ( .D(n708), .CLK(clk), .Q(\mem[18][18] ) );
  DFFX1 \mem_reg[18][17]  ( .D(n707), .CLK(clk), .Q(\mem[18][17] ) );
  DFFX1 \mem_reg[18][16]  ( .D(n706), .CLK(clk), .Q(\mem[18][16] ) );
  DFFX1 \mem_reg[18][15]  ( .D(n705), .CLK(clk), .Q(\mem[18][15] ) );
  DFFX1 \mem_reg[18][14]  ( .D(n704), .CLK(clk), .Q(\mem[18][14] ) );
  DFFX1 \mem_reg[18][13]  ( .D(n703), .CLK(clk), .Q(\mem[18][13] ) );
  DFFX1 \mem_reg[18][12]  ( .D(n702), .CLK(clk), .Q(\mem[18][12] ) );
  DFFX1 \mem_reg[18][11]  ( .D(n701), .CLK(clk), .Q(\mem[18][11] ) );
  DFFX1 \mem_reg[18][10]  ( .D(n700), .CLK(clk), .Q(\mem[18][10] ) );
  DFFX1 \mem_reg[18][9]  ( .D(n699), .CLK(clk), .Q(\mem[18][9] ) );
  DFFX1 \mem_reg[18][8]  ( .D(n698), .CLK(clk), .Q(\mem[18][8] ) );
  DFFX1 \mem_reg[18][7]  ( .D(n697), .CLK(clk), .Q(\mem[18][7] ) );
  DFFX1 \mem_reg[18][6]  ( .D(n696), .CLK(clk), .Q(\mem[18][6] ) );
  DFFX1 \mem_reg[18][5]  ( .D(n695), .CLK(clk), .Q(\mem[18][5] ) );
  DFFX1 \mem_reg[18][4]  ( .D(n694), .CLK(clk), .Q(\mem[18][4] ) );
  DFFX1 \mem_reg[18][3]  ( .D(n693), .CLK(clk), .Q(\mem[18][3] ) );
  DFFX1 \mem_reg[18][2]  ( .D(n692), .CLK(clk), .Q(\mem[18][2] ) );
  DFFX1 \mem_reg[18][1]  ( .D(n691), .CLK(clk), .Q(\mem[18][1] ) );
  DFFX1 \mem_reg[18][0]  ( .D(n690), .CLK(clk), .Q(\mem[18][0] ) );
  DFFX1 \mem_reg[17][31]  ( .D(n689), .CLK(clk), .Q(\mem[17][31] ) );
  DFFX1 \mem_reg[17][30]  ( .D(n688), .CLK(clk), .Q(\mem[17][30] ) );
  DFFX1 \mem_reg[17][29]  ( .D(n687), .CLK(clk), .Q(\mem[17][29] ) );
  DFFX1 \mem_reg[17][28]  ( .D(n686), .CLK(clk), .Q(\mem[17][28] ) );
  DFFX1 \mem_reg[17][27]  ( .D(n685), .CLK(clk), .Q(\mem[17][27] ) );
  DFFX1 \mem_reg[17][26]  ( .D(n684), .CLK(clk), .Q(\mem[17][26] ) );
  DFFX1 \mem_reg[17][25]  ( .D(n683), .CLK(clk), .Q(\mem[17][25] ) );
  DFFX1 \mem_reg[17][24]  ( .D(n682), .CLK(clk), .Q(\mem[17][24] ) );
  DFFX1 \mem_reg[17][23]  ( .D(n681), .CLK(clk), .Q(\mem[17][23] ) );
  DFFX1 \mem_reg[17][22]  ( .D(n680), .CLK(clk), .Q(\mem[17][22] ) );
  DFFX1 \mem_reg[17][21]  ( .D(n679), .CLK(clk), .Q(\mem[17][21] ) );
  DFFX1 \mem_reg[17][20]  ( .D(n678), .CLK(clk), .Q(\mem[17][20] ) );
  DFFX1 \mem_reg[17][19]  ( .D(n677), .CLK(clk), .Q(\mem[17][19] ) );
  DFFX1 \mem_reg[17][18]  ( .D(n676), .CLK(clk), .Q(\mem[17][18] ) );
  DFFX1 \mem_reg[17][17]  ( .D(n675), .CLK(clk), .Q(\mem[17][17] ) );
  DFFX1 \mem_reg[17][16]  ( .D(n674), .CLK(clk), .Q(\mem[17][16] ) );
  DFFX1 \mem_reg[17][15]  ( .D(n673), .CLK(clk), .Q(\mem[17][15] ) );
  DFFX1 \mem_reg[17][14]  ( .D(n672), .CLK(clk), .Q(\mem[17][14] ) );
  DFFX1 \mem_reg[17][13]  ( .D(n671), .CLK(clk), .Q(\mem[17][13] ) );
  DFFX1 \mem_reg[17][12]  ( .D(n670), .CLK(clk), .Q(\mem[17][12] ) );
  DFFX1 \mem_reg[17][11]  ( .D(n669), .CLK(clk), .Q(\mem[17][11] ) );
  DFFX1 \mem_reg[17][10]  ( .D(n668), .CLK(clk), .Q(\mem[17][10] ) );
  DFFX1 \mem_reg[17][9]  ( .D(n667), .CLK(clk), .Q(\mem[17][9] ) );
  DFFX1 \mem_reg[17][8]  ( .D(n666), .CLK(clk), .Q(\mem[17][8] ) );
  DFFX1 \mem_reg[17][7]  ( .D(n665), .CLK(clk), .Q(\mem[17][7] ) );
  DFFX1 \mem_reg[17][6]  ( .D(n664), .CLK(clk), .Q(\mem[17][6] ) );
  DFFX1 \mem_reg[17][5]  ( .D(n663), .CLK(clk), .Q(\mem[17][5] ) );
  DFFX1 \mem_reg[17][4]  ( .D(n662), .CLK(clk), .Q(\mem[17][4] ) );
  DFFX1 \mem_reg[17][3]  ( .D(n661), .CLK(clk), .Q(\mem[17][3] ) );
  DFFX1 \mem_reg[17][2]  ( .D(n660), .CLK(clk), .Q(\mem[17][2] ) );
  DFFX1 \mem_reg[17][1]  ( .D(n659), .CLK(clk), .Q(\mem[17][1] ) );
  DFFX1 \mem_reg[17][0]  ( .D(n658), .CLK(clk), .Q(\mem[17][0] ) );
  DFFX1 \mem_reg[16][31]  ( .D(n657), .CLK(clk), .Q(\mem[16][31] ) );
  DFFX1 \mem_reg[16][30]  ( .D(n656), .CLK(clk), .Q(\mem[16][30] ) );
  DFFX1 \mem_reg[16][29]  ( .D(n655), .CLK(clk), .Q(\mem[16][29] ) );
  DFFX1 \mem_reg[16][28]  ( .D(n654), .CLK(clk), .Q(\mem[16][28] ) );
  DFFX1 \mem_reg[16][27]  ( .D(n653), .CLK(clk), .Q(\mem[16][27] ) );
  DFFX1 \mem_reg[16][26]  ( .D(n652), .CLK(clk), .Q(\mem[16][26] ) );
  DFFX1 \mem_reg[16][25]  ( .D(n651), .CLK(clk), .Q(\mem[16][25] ) );
  DFFX1 \mem_reg[16][24]  ( .D(n650), .CLK(clk), .Q(\mem[16][24] ) );
  DFFX1 \mem_reg[16][23]  ( .D(n649), .CLK(clk), .Q(\mem[16][23] ) );
  DFFX1 \mem_reg[16][22]  ( .D(n648), .CLK(clk), .Q(\mem[16][22] ) );
  DFFX1 \mem_reg[16][21]  ( .D(n647), .CLK(clk), .Q(\mem[16][21] ) );
  DFFX1 \mem_reg[16][20]  ( .D(n646), .CLK(clk), .Q(\mem[16][20] ) );
  DFFX1 \mem_reg[16][19]  ( .D(n645), .CLK(clk), .Q(\mem[16][19] ) );
  DFFX1 \mem_reg[16][18]  ( .D(n644), .CLK(clk), .Q(\mem[16][18] ) );
  DFFX1 \mem_reg[16][17]  ( .D(n643), .CLK(clk), .Q(\mem[16][17] ) );
  DFFX1 \mem_reg[16][16]  ( .D(n642), .CLK(clk), .Q(\mem[16][16] ) );
  DFFX1 \mem_reg[16][15]  ( .D(n641), .CLK(clk), .Q(\mem[16][15] ) );
  DFFX1 \mem_reg[16][14]  ( .D(n640), .CLK(clk), .Q(\mem[16][14] ) );
  DFFX1 \mem_reg[16][13]  ( .D(n639), .CLK(clk), .Q(\mem[16][13] ) );
  DFFX1 \mem_reg[16][12]  ( .D(n638), .CLK(clk), .Q(\mem[16][12] ) );
  DFFX1 \mem_reg[16][11]  ( .D(n637), .CLK(clk), .Q(\mem[16][11] ) );
  DFFX1 \mem_reg[16][10]  ( .D(n636), .CLK(clk), .Q(\mem[16][10] ) );
  DFFX1 \mem_reg[16][9]  ( .D(n635), .CLK(clk), .Q(\mem[16][9] ) );
  DFFX1 \mem_reg[16][8]  ( .D(n634), .CLK(clk), .Q(\mem[16][8] ) );
  DFFX1 \mem_reg[16][7]  ( .D(n633), .CLK(clk), .Q(\mem[16][7] ) );
  DFFX1 \mem_reg[16][6]  ( .D(n632), .CLK(clk), .Q(\mem[16][6] ) );
  DFFX1 \mem_reg[16][5]  ( .D(n631), .CLK(clk), .Q(\mem[16][5] ) );
  DFFX1 \mem_reg[16][4]  ( .D(n630), .CLK(clk), .Q(\mem[16][4] ) );
  DFFX1 \mem_reg[16][3]  ( .D(n629), .CLK(clk), .Q(\mem[16][3] ) );
  DFFX1 \mem_reg[16][2]  ( .D(n628), .CLK(clk), .Q(\mem[16][2] ) );
  DFFX1 \mem_reg[16][1]  ( .D(n627), .CLK(clk), .Q(\mem[16][1] ) );
  DFFX1 \mem_reg[16][0]  ( .D(n626), .CLK(clk), .Q(\mem[16][0] ) );
  DFFX1 \mem_reg[15][31]  ( .D(n625), .CLK(clk), .Q(\mem[15][31] ) );
  DFFX1 \mem_reg[15][30]  ( .D(n624), .CLK(clk), .Q(\mem[15][30] ) );
  DFFX1 \mem_reg[15][29]  ( .D(n623), .CLK(clk), .Q(\mem[15][29] ) );
  DFFX1 \mem_reg[15][28]  ( .D(n622), .CLK(clk), .Q(\mem[15][28] ) );
  DFFX1 \mem_reg[15][27]  ( .D(n621), .CLK(clk), .Q(\mem[15][27] ) );
  DFFX1 \mem_reg[15][26]  ( .D(n620), .CLK(clk), .Q(\mem[15][26] ) );
  DFFX1 \mem_reg[15][25]  ( .D(n619), .CLK(clk), .Q(\mem[15][25] ) );
  DFFX1 \mem_reg[15][24]  ( .D(n618), .CLK(clk), .Q(\mem[15][24] ) );
  DFFX1 \mem_reg[15][23]  ( .D(n617), .CLK(clk), .Q(\mem[15][23] ) );
  DFFX1 \mem_reg[15][22]  ( .D(n616), .CLK(clk), .Q(\mem[15][22] ) );
  DFFX1 \mem_reg[15][21]  ( .D(n615), .CLK(clk), .Q(\mem[15][21] ) );
  DFFX1 \mem_reg[15][20]  ( .D(n614), .CLK(clk), .Q(\mem[15][20] ) );
  DFFX1 \mem_reg[15][19]  ( .D(n613), .CLK(clk), .Q(\mem[15][19] ) );
  DFFX1 \mem_reg[15][18]  ( .D(n612), .CLK(clk), .Q(\mem[15][18] ) );
  DFFX1 \mem_reg[15][17]  ( .D(n611), .CLK(clk), .Q(\mem[15][17] ) );
  DFFX1 \mem_reg[15][16]  ( .D(n610), .CLK(clk), .Q(\mem[15][16] ) );
  DFFX1 \mem_reg[15][15]  ( .D(n609), .CLK(clk), .Q(\mem[15][15] ) );
  DFFX1 \mem_reg[15][14]  ( .D(n608), .CLK(clk), .Q(\mem[15][14] ) );
  DFFX1 \mem_reg[15][13]  ( .D(n607), .CLK(clk), .Q(\mem[15][13] ) );
  DFFX1 \mem_reg[15][12]  ( .D(n606), .CLK(clk), .Q(\mem[15][12] ) );
  DFFX1 \mem_reg[15][11]  ( .D(n605), .CLK(clk), .Q(\mem[15][11] ) );
  DFFX1 \mem_reg[15][10]  ( .D(n604), .CLK(clk), .Q(\mem[15][10] ) );
  DFFX1 \mem_reg[15][9]  ( .D(n603), .CLK(clk), .Q(\mem[15][9] ) );
  DFFX1 \mem_reg[15][8]  ( .D(n602), .CLK(clk), .Q(\mem[15][8] ) );
  DFFX1 \mem_reg[15][7]  ( .D(n601), .CLK(clk), .Q(\mem[15][7] ) );
  DFFX1 \mem_reg[15][6]  ( .D(n600), .CLK(clk), .Q(\mem[15][6] ) );
  DFFX1 \mem_reg[15][5]  ( .D(n599), .CLK(clk), .Q(\mem[15][5] ) );
  DFFX1 \mem_reg[15][4]  ( .D(n598), .CLK(clk), .Q(\mem[15][4] ) );
  DFFX1 \mem_reg[15][3]  ( .D(n597), .CLK(clk), .Q(\mem[15][3] ) );
  DFFX1 \mem_reg[15][2]  ( .D(n596), .CLK(clk), .Q(\mem[15][2] ) );
  DFFX1 \mem_reg[15][1]  ( .D(n595), .CLK(clk), .Q(\mem[15][1] ) );
  DFFX1 \mem_reg[15][0]  ( .D(n594), .CLK(clk), .Q(\mem[15][0] ) );
  DFFX1 \mem_reg[14][31]  ( .D(n593), .CLK(clk), .Q(\mem[14][31] ) );
  DFFX1 \mem_reg[14][30]  ( .D(n592), .CLK(clk), .Q(\mem[14][30] ) );
  DFFX1 \mem_reg[14][29]  ( .D(n591), .CLK(clk), .Q(\mem[14][29] ) );
  DFFX1 \mem_reg[14][28]  ( .D(n590), .CLK(clk), .Q(\mem[14][28] ) );
  DFFX1 \mem_reg[14][27]  ( .D(n589), .CLK(clk), .Q(\mem[14][27] ) );
  DFFX1 \mem_reg[14][26]  ( .D(n588), .CLK(clk), .Q(\mem[14][26] ) );
  DFFX1 \mem_reg[14][25]  ( .D(n587), .CLK(clk), .Q(\mem[14][25] ) );
  DFFX1 \mem_reg[14][24]  ( .D(n586), .CLK(clk), .Q(\mem[14][24] ) );
  DFFX1 \mem_reg[14][23]  ( .D(n585), .CLK(clk), .Q(\mem[14][23] ) );
  DFFX1 \mem_reg[14][22]  ( .D(n584), .CLK(clk), .Q(\mem[14][22] ) );
  DFFX1 \mem_reg[14][21]  ( .D(n583), .CLK(clk), .Q(\mem[14][21] ) );
  DFFX1 \mem_reg[14][20]  ( .D(n582), .CLK(clk), .Q(\mem[14][20] ) );
  DFFX1 \mem_reg[14][19]  ( .D(n581), .CLK(clk), .Q(\mem[14][19] ) );
  DFFX1 \mem_reg[14][18]  ( .D(n580), .CLK(clk), .Q(\mem[14][18] ) );
  DFFX1 \mem_reg[14][17]  ( .D(n579), .CLK(clk), .Q(\mem[14][17] ) );
  DFFX1 \mem_reg[14][16]  ( .D(n578), .CLK(clk), .Q(\mem[14][16] ) );
  DFFX1 \mem_reg[14][15]  ( .D(n577), .CLK(clk), .Q(\mem[14][15] ) );
  DFFX1 \mem_reg[14][14]  ( .D(n576), .CLK(clk), .Q(\mem[14][14] ) );
  DFFX1 \mem_reg[14][13]  ( .D(n575), .CLK(clk), .Q(\mem[14][13] ) );
  DFFX1 \mem_reg[14][12]  ( .D(n574), .CLK(clk), .Q(\mem[14][12] ) );
  DFFX1 \mem_reg[14][11]  ( .D(n573), .CLK(clk), .Q(\mem[14][11] ) );
  DFFX1 \mem_reg[14][10]  ( .D(n572), .CLK(clk), .Q(\mem[14][10] ) );
  DFFX1 \mem_reg[14][9]  ( .D(n571), .CLK(clk), .Q(\mem[14][9] ) );
  DFFX1 \mem_reg[14][8]  ( .D(n570), .CLK(clk), .Q(\mem[14][8] ) );
  DFFX1 \mem_reg[14][7]  ( .D(n569), .CLK(clk), .Q(\mem[14][7] ) );
  DFFX1 \mem_reg[14][6]  ( .D(n568), .CLK(clk), .Q(\mem[14][6] ) );
  DFFX1 \mem_reg[14][5]  ( .D(n567), .CLK(clk), .Q(\mem[14][5] ) );
  DFFX1 \mem_reg[14][4]  ( .D(n566), .CLK(clk), .Q(\mem[14][4] ) );
  DFFX1 \mem_reg[14][3]  ( .D(n565), .CLK(clk), .Q(\mem[14][3] ) );
  DFFX1 \mem_reg[14][2]  ( .D(n564), .CLK(clk), .Q(\mem[14][2] ) );
  DFFX1 \mem_reg[14][1]  ( .D(n563), .CLK(clk), .Q(\mem[14][1] ) );
  DFFX1 \mem_reg[14][0]  ( .D(n562), .CLK(clk), .Q(\mem[14][0] ) );
  DFFX1 \mem_reg[13][31]  ( .D(n561), .CLK(clk), .Q(\mem[13][31] ) );
  DFFX1 \mem_reg[13][30]  ( .D(n560), .CLK(clk), .Q(\mem[13][30] ) );
  DFFX1 \mem_reg[13][29]  ( .D(n559), .CLK(clk), .Q(\mem[13][29] ) );
  DFFX1 \mem_reg[13][28]  ( .D(n558), .CLK(clk), .Q(\mem[13][28] ) );
  DFFX1 \mem_reg[13][27]  ( .D(n557), .CLK(clk), .Q(\mem[13][27] ) );
  DFFX1 \mem_reg[13][26]  ( .D(n556), .CLK(clk), .Q(\mem[13][26] ) );
  DFFX1 \mem_reg[13][25]  ( .D(n555), .CLK(clk), .Q(\mem[13][25] ) );
  DFFX1 \mem_reg[13][24]  ( .D(n554), .CLK(clk), .Q(\mem[13][24] ) );
  DFFX1 \mem_reg[13][23]  ( .D(n553), .CLK(clk), .Q(\mem[13][23] ) );
  DFFX1 \mem_reg[13][22]  ( .D(n552), .CLK(clk), .Q(\mem[13][22] ) );
  DFFX1 \mem_reg[13][21]  ( .D(n551), .CLK(clk), .Q(\mem[13][21] ) );
  DFFX1 \mem_reg[13][20]  ( .D(n550), .CLK(clk), .Q(\mem[13][20] ) );
  DFFX1 \mem_reg[13][19]  ( .D(n549), .CLK(clk), .Q(\mem[13][19] ) );
  DFFX1 \mem_reg[13][18]  ( .D(n548), .CLK(clk), .Q(\mem[13][18] ) );
  DFFX1 \mem_reg[13][17]  ( .D(n547), .CLK(clk), .Q(\mem[13][17] ) );
  DFFX1 \mem_reg[13][16]  ( .D(n546), .CLK(clk), .Q(\mem[13][16] ) );
  DFFX1 \mem_reg[13][15]  ( .D(n545), .CLK(clk), .Q(\mem[13][15] ) );
  DFFX1 \mem_reg[13][14]  ( .D(n544), .CLK(clk), .Q(\mem[13][14] ) );
  DFFX1 \mem_reg[13][13]  ( .D(n543), .CLK(clk), .Q(\mem[13][13] ) );
  DFFX1 \mem_reg[13][12]  ( .D(n542), .CLK(clk), .Q(\mem[13][12] ) );
  DFFX1 \mem_reg[13][11]  ( .D(n541), .CLK(clk), .Q(\mem[13][11] ) );
  DFFX1 \mem_reg[13][10]  ( .D(n540), .CLK(clk), .Q(\mem[13][10] ) );
  DFFX1 \mem_reg[13][9]  ( .D(n539), .CLK(clk), .Q(\mem[13][9] ) );
  DFFX1 \mem_reg[13][8]  ( .D(n538), .CLK(clk), .Q(\mem[13][8] ) );
  DFFX1 \mem_reg[13][7]  ( .D(n537), .CLK(clk), .Q(\mem[13][7] ) );
  DFFX1 \mem_reg[13][6]  ( .D(n536), .CLK(clk), .Q(\mem[13][6] ) );
  DFFX1 \mem_reg[13][5]  ( .D(n535), .CLK(clk), .Q(\mem[13][5] ) );
  DFFX1 \mem_reg[13][4]  ( .D(n534), .CLK(clk), .Q(\mem[13][4] ) );
  DFFX1 \mem_reg[13][3]  ( .D(n533), .CLK(clk), .Q(\mem[13][3] ) );
  DFFX1 \mem_reg[13][2]  ( .D(n532), .CLK(clk), .Q(\mem[13][2] ) );
  DFFX1 \mem_reg[13][1]  ( .D(n531), .CLK(clk), .Q(\mem[13][1] ) );
  DFFX1 \mem_reg[13][0]  ( .D(n530), .CLK(clk), .Q(\mem[13][0] ) );
  DFFX1 \mem_reg[12][31]  ( .D(n529), .CLK(clk), .Q(\mem[12][31] ) );
  DFFX1 \mem_reg[12][30]  ( .D(n528), .CLK(clk), .Q(\mem[12][30] ) );
  DFFX1 \mem_reg[12][29]  ( .D(n527), .CLK(clk), .Q(\mem[12][29] ) );
  DFFX1 \mem_reg[12][28]  ( .D(n526), .CLK(clk), .Q(\mem[12][28] ) );
  DFFX1 \mem_reg[12][27]  ( .D(n525), .CLK(clk), .Q(\mem[12][27] ) );
  DFFX1 \mem_reg[12][26]  ( .D(n524), .CLK(clk), .Q(\mem[12][26] ) );
  DFFX1 \mem_reg[12][25]  ( .D(n523), .CLK(clk), .Q(\mem[12][25] ) );
  DFFX1 \mem_reg[12][24]  ( .D(n522), .CLK(clk), .Q(\mem[12][24] ) );
  DFFX1 \mem_reg[12][23]  ( .D(n521), .CLK(clk), .Q(\mem[12][23] ) );
  DFFX1 \mem_reg[12][22]  ( .D(n520), .CLK(clk), .Q(\mem[12][22] ) );
  DFFX1 \mem_reg[12][21]  ( .D(n519), .CLK(clk), .Q(\mem[12][21] ) );
  DFFX1 \mem_reg[12][20]  ( .D(n518), .CLK(clk), .Q(\mem[12][20] ) );
  DFFX1 \mem_reg[12][19]  ( .D(n517), .CLK(clk), .Q(\mem[12][19] ) );
  DFFX1 \mem_reg[12][18]  ( .D(n516), .CLK(clk), .Q(\mem[12][18] ) );
  DFFX1 \mem_reg[12][17]  ( .D(n515), .CLK(clk), .Q(\mem[12][17] ) );
  DFFX1 \mem_reg[12][16]  ( .D(n514), .CLK(clk), .Q(\mem[12][16] ) );
  DFFX1 \mem_reg[12][15]  ( .D(n513), .CLK(clk), .Q(\mem[12][15] ) );
  DFFX1 \mem_reg[12][14]  ( .D(n512), .CLK(clk), .Q(\mem[12][14] ) );
  DFFX1 \mem_reg[12][13]  ( .D(n511), .CLK(clk), .Q(\mem[12][13] ) );
  DFFX1 \mem_reg[12][12]  ( .D(n510), .CLK(clk), .Q(\mem[12][12] ) );
  DFFX1 \mem_reg[12][11]  ( .D(n509), .CLK(clk), .Q(\mem[12][11] ) );
  DFFX1 \mem_reg[12][10]  ( .D(n508), .CLK(clk), .Q(\mem[12][10] ) );
  DFFX1 \mem_reg[12][9]  ( .D(n507), .CLK(clk), .Q(\mem[12][9] ) );
  DFFX1 \mem_reg[12][8]  ( .D(n506), .CLK(clk), .Q(\mem[12][8] ) );
  DFFX1 \mem_reg[12][7]  ( .D(n505), .CLK(clk), .Q(\mem[12][7] ) );
  DFFX1 \mem_reg[12][6]  ( .D(n504), .CLK(clk), .Q(\mem[12][6] ) );
  DFFX1 \mem_reg[12][5]  ( .D(n503), .CLK(clk), .Q(\mem[12][5] ) );
  DFFX1 \mem_reg[12][4]  ( .D(n502), .CLK(clk), .Q(\mem[12][4] ) );
  DFFX1 \mem_reg[12][3]  ( .D(n501), .CLK(clk), .Q(\mem[12][3] ) );
  DFFX1 \mem_reg[12][2]  ( .D(n500), .CLK(clk), .Q(\mem[12][2] ) );
  DFFX1 \mem_reg[12][1]  ( .D(n499), .CLK(clk), .Q(\mem[12][1] ) );
  DFFX1 \mem_reg[12][0]  ( .D(n498), .CLK(clk), .Q(\mem[12][0] ) );
  DFFX1 \mem_reg[11][31]  ( .D(n497), .CLK(clk), .Q(\mem[11][31] ) );
  DFFX1 \mem_reg[11][30]  ( .D(n496), .CLK(clk), .Q(\mem[11][30] ) );
  DFFX1 \mem_reg[11][29]  ( .D(n495), .CLK(clk), .Q(\mem[11][29] ) );
  DFFX1 \mem_reg[11][28]  ( .D(n494), .CLK(clk), .Q(\mem[11][28] ) );
  DFFX1 \mem_reg[11][27]  ( .D(n493), .CLK(clk), .Q(\mem[11][27] ) );
  DFFX1 \mem_reg[11][26]  ( .D(n492), .CLK(clk), .Q(\mem[11][26] ) );
  DFFX1 \mem_reg[11][25]  ( .D(n491), .CLK(clk), .Q(\mem[11][25] ) );
  DFFX1 \mem_reg[11][24]  ( .D(n490), .CLK(clk), .Q(\mem[11][24] ) );
  DFFX1 \mem_reg[11][23]  ( .D(n489), .CLK(clk), .Q(\mem[11][23] ) );
  DFFX1 \mem_reg[11][22]  ( .D(n488), .CLK(clk), .Q(\mem[11][22] ) );
  DFFX1 \mem_reg[11][21]  ( .D(n487), .CLK(clk), .Q(\mem[11][21] ) );
  DFFX1 \mem_reg[11][20]  ( .D(n486), .CLK(clk), .Q(\mem[11][20] ) );
  DFFX1 \mem_reg[11][19]  ( .D(n485), .CLK(clk), .Q(\mem[11][19] ) );
  DFFX1 \mem_reg[11][18]  ( .D(n484), .CLK(clk), .Q(\mem[11][18] ) );
  DFFX1 \mem_reg[11][17]  ( .D(n483), .CLK(clk), .Q(\mem[11][17] ) );
  DFFX1 \mem_reg[11][16]  ( .D(n482), .CLK(clk), .Q(\mem[11][16] ) );
  DFFX1 \mem_reg[11][15]  ( .D(n481), .CLK(clk), .Q(\mem[11][15] ) );
  DFFX1 \mem_reg[11][14]  ( .D(n480), .CLK(clk), .Q(\mem[11][14] ) );
  DFFX1 \mem_reg[11][13]  ( .D(n479), .CLK(clk), .Q(\mem[11][13] ) );
  DFFX1 \mem_reg[11][12]  ( .D(n478), .CLK(clk), .Q(\mem[11][12] ) );
  DFFX1 \mem_reg[11][11]  ( .D(n477), .CLK(clk), .Q(\mem[11][11] ) );
  DFFX1 \mem_reg[11][10]  ( .D(n476), .CLK(clk), .Q(\mem[11][10] ) );
  DFFX1 \mem_reg[11][9]  ( .D(n475), .CLK(clk), .Q(\mem[11][9] ) );
  DFFX1 \mem_reg[11][8]  ( .D(n474), .CLK(clk), .Q(\mem[11][8] ) );
  DFFX1 \mem_reg[11][7]  ( .D(n473), .CLK(clk), .Q(\mem[11][7] ) );
  DFFX1 \mem_reg[11][6]  ( .D(n472), .CLK(clk), .Q(\mem[11][6] ) );
  DFFX1 \mem_reg[11][5]  ( .D(n471), .CLK(clk), .Q(\mem[11][5] ) );
  DFFX1 \mem_reg[11][4]  ( .D(n470), .CLK(clk), .Q(\mem[11][4] ) );
  DFFX1 \mem_reg[11][3]  ( .D(n469), .CLK(clk), .Q(\mem[11][3] ) );
  DFFX1 \mem_reg[11][2]  ( .D(n468), .CLK(clk), .Q(\mem[11][2] ) );
  DFFX1 \mem_reg[11][1]  ( .D(n467), .CLK(clk), .Q(\mem[11][1] ) );
  DFFX1 \mem_reg[11][0]  ( .D(n466), .CLK(clk), .Q(\mem[11][0] ) );
  DFFX1 \mem_reg[10][31]  ( .D(n465), .CLK(clk), .Q(\mem[10][31] ) );
  DFFX1 \mem_reg[10][30]  ( .D(n464), .CLK(clk), .Q(\mem[10][30] ) );
  DFFX1 \mem_reg[10][29]  ( .D(n463), .CLK(clk), .Q(\mem[10][29] ) );
  DFFX1 \mem_reg[10][28]  ( .D(n462), .CLK(clk), .Q(\mem[10][28] ) );
  DFFX1 \mem_reg[10][27]  ( .D(n461), .CLK(clk), .Q(\mem[10][27] ) );
  DFFX1 \mem_reg[10][26]  ( .D(n460), .CLK(clk), .Q(\mem[10][26] ) );
  DFFX1 \mem_reg[10][25]  ( .D(n459), .CLK(clk), .Q(\mem[10][25] ) );
  DFFX1 \mem_reg[10][24]  ( .D(n458), .CLK(clk), .Q(\mem[10][24] ) );
  DFFX1 \mem_reg[10][23]  ( .D(n457), .CLK(clk), .Q(\mem[10][23] ) );
  DFFX1 \mem_reg[10][22]  ( .D(n456), .CLK(clk), .Q(\mem[10][22] ) );
  DFFX1 \mem_reg[10][21]  ( .D(n455), .CLK(clk), .Q(\mem[10][21] ) );
  DFFX1 \mem_reg[10][20]  ( .D(n454), .CLK(clk), .Q(\mem[10][20] ) );
  DFFX1 \mem_reg[10][19]  ( .D(n453), .CLK(clk), .Q(\mem[10][19] ) );
  DFFX1 \mem_reg[10][18]  ( .D(n452), .CLK(clk), .Q(\mem[10][18] ) );
  DFFX1 \mem_reg[10][17]  ( .D(n451), .CLK(clk), .Q(\mem[10][17] ) );
  DFFX1 \mem_reg[10][16]  ( .D(n450), .CLK(clk), .Q(\mem[10][16] ) );
  DFFX1 \mem_reg[10][15]  ( .D(n449), .CLK(clk), .Q(\mem[10][15] ) );
  DFFX1 \mem_reg[10][14]  ( .D(n448), .CLK(clk), .Q(\mem[10][14] ) );
  DFFX1 \mem_reg[10][13]  ( .D(n447), .CLK(clk), .Q(\mem[10][13] ) );
  DFFX1 \mem_reg[10][12]  ( .D(n446), .CLK(clk), .Q(\mem[10][12] ) );
  DFFX1 \mem_reg[10][11]  ( .D(n445), .CLK(clk), .Q(\mem[10][11] ) );
  DFFX1 \mem_reg[10][10]  ( .D(n444), .CLK(clk), .Q(\mem[10][10] ) );
  DFFX1 \mem_reg[10][9]  ( .D(n443), .CLK(clk), .Q(\mem[10][9] ) );
  DFFX1 \mem_reg[10][8]  ( .D(n442), .CLK(clk), .Q(\mem[10][8] ) );
  DFFX1 \mem_reg[10][7]  ( .D(n441), .CLK(clk), .Q(\mem[10][7] ) );
  DFFX1 \mem_reg[10][6]  ( .D(n440), .CLK(clk), .Q(\mem[10][6] ) );
  DFFX1 \mem_reg[10][5]  ( .D(n439), .CLK(clk), .Q(\mem[10][5] ) );
  DFFX1 \mem_reg[10][4]  ( .D(n438), .CLK(clk), .Q(\mem[10][4] ) );
  DFFX1 \mem_reg[10][3]  ( .D(n437), .CLK(clk), .Q(\mem[10][3] ) );
  DFFX1 \mem_reg[10][2]  ( .D(n436), .CLK(clk), .Q(\mem[10][2] ) );
  DFFX1 \mem_reg[10][1]  ( .D(n435), .CLK(clk), .Q(\mem[10][1] ) );
  DFFX1 \mem_reg[10][0]  ( .D(n434), .CLK(clk), .Q(\mem[10][0] ) );
  DFFX1 \mem_reg[9][31]  ( .D(n433), .CLK(clk), .Q(\mem[9][31] ) );
  DFFX1 \mem_reg[9][30]  ( .D(n432), .CLK(clk), .Q(\mem[9][30] ) );
  DFFX1 \mem_reg[9][29]  ( .D(n431), .CLK(clk), .Q(\mem[9][29] ) );
  DFFX1 \mem_reg[9][28]  ( .D(n430), .CLK(clk), .Q(\mem[9][28] ) );
  DFFX1 \mem_reg[9][27]  ( .D(n429), .CLK(clk), .Q(\mem[9][27] ) );
  DFFX1 \mem_reg[9][26]  ( .D(n428), .CLK(clk), .Q(\mem[9][26] ) );
  DFFX1 \mem_reg[9][25]  ( .D(n427), .CLK(clk), .Q(\mem[9][25] ) );
  DFFX1 \mem_reg[9][24]  ( .D(n426), .CLK(clk), .Q(\mem[9][24] ) );
  DFFX1 \mem_reg[9][23]  ( .D(n425), .CLK(clk), .Q(\mem[9][23] ) );
  DFFX1 \mem_reg[9][22]  ( .D(n424), .CLK(clk), .Q(\mem[9][22] ) );
  DFFX1 \mem_reg[9][21]  ( .D(n423), .CLK(clk), .Q(\mem[9][21] ) );
  DFFX1 \mem_reg[9][20]  ( .D(n422), .CLK(clk), .Q(\mem[9][20] ) );
  DFFX1 \mem_reg[9][19]  ( .D(n421), .CLK(clk), .Q(\mem[9][19] ) );
  DFFX1 \mem_reg[9][18]  ( .D(n420), .CLK(clk), .Q(\mem[9][18] ) );
  DFFX1 \mem_reg[9][17]  ( .D(n419), .CLK(clk), .Q(\mem[9][17] ) );
  DFFX1 \mem_reg[9][16]  ( .D(n418), .CLK(clk), .Q(\mem[9][16] ) );
  DFFX1 \mem_reg[9][15]  ( .D(n417), .CLK(clk), .Q(\mem[9][15] ) );
  DFFX1 \mem_reg[9][14]  ( .D(n416), .CLK(clk), .Q(\mem[9][14] ) );
  DFFX1 \mem_reg[9][13]  ( .D(n415), .CLK(clk), .Q(\mem[9][13] ) );
  DFFX1 \mem_reg[9][12]  ( .D(n414), .CLK(clk), .Q(\mem[9][12] ) );
  DFFX1 \mem_reg[9][11]  ( .D(n413), .CLK(clk), .Q(\mem[9][11] ) );
  DFFX1 \mem_reg[9][10]  ( .D(n412), .CLK(clk), .Q(\mem[9][10] ) );
  DFFX1 \mem_reg[9][9]  ( .D(n411), .CLK(clk), .Q(\mem[9][9] ) );
  DFFX1 \mem_reg[9][8]  ( .D(n410), .CLK(clk), .Q(\mem[9][8] ) );
  DFFX1 \mem_reg[9][7]  ( .D(n409), .CLK(clk), .Q(\mem[9][7] ) );
  DFFX1 \mem_reg[9][6]  ( .D(n408), .CLK(clk), .Q(\mem[9][6] ) );
  DFFX1 \mem_reg[9][5]  ( .D(n407), .CLK(clk), .Q(\mem[9][5] ) );
  DFFX1 \mem_reg[9][4]  ( .D(n406), .CLK(clk), .Q(\mem[9][4] ) );
  DFFX1 \mem_reg[9][3]  ( .D(n405), .CLK(clk), .Q(\mem[9][3] ) );
  DFFX1 \mem_reg[9][2]  ( .D(n404), .CLK(clk), .Q(\mem[9][2] ) );
  DFFX1 \mem_reg[9][1]  ( .D(n403), .CLK(clk), .Q(\mem[9][1] ) );
  DFFX1 \mem_reg[9][0]  ( .D(n402), .CLK(clk), .Q(\mem[9][0] ) );
  DFFX1 \mem_reg[8][31]  ( .D(n401), .CLK(clk), .Q(\mem[8][31] ) );
  DFFX1 \mem_reg[8][30]  ( .D(n400), .CLK(clk), .Q(\mem[8][30] ) );
  DFFX1 \mem_reg[8][29]  ( .D(n399), .CLK(clk), .Q(\mem[8][29] ) );
  DFFX1 \mem_reg[8][28]  ( .D(n398), .CLK(clk), .Q(\mem[8][28] ) );
  DFFX1 \mem_reg[8][27]  ( .D(n397), .CLK(clk), .Q(\mem[8][27] ) );
  DFFX1 \mem_reg[8][26]  ( .D(n396), .CLK(clk), .Q(\mem[8][26] ) );
  DFFX1 \mem_reg[8][25]  ( .D(n395), .CLK(clk), .Q(\mem[8][25] ) );
  DFFX1 \mem_reg[8][24]  ( .D(n394), .CLK(clk), .Q(\mem[8][24] ) );
  DFFX1 \mem_reg[8][23]  ( .D(n393), .CLK(clk), .Q(\mem[8][23] ) );
  DFFX1 \mem_reg[8][22]  ( .D(n392), .CLK(clk), .Q(\mem[8][22] ) );
  DFFX1 \mem_reg[8][21]  ( .D(n391), .CLK(clk), .Q(\mem[8][21] ) );
  DFFX1 \mem_reg[8][20]  ( .D(n390), .CLK(clk), .Q(\mem[8][20] ) );
  DFFX1 \mem_reg[8][19]  ( .D(n389), .CLK(clk), .Q(\mem[8][19] ) );
  DFFX1 \mem_reg[8][18]  ( .D(n388), .CLK(clk), .Q(\mem[8][18] ) );
  DFFX1 \mem_reg[8][17]  ( .D(n387), .CLK(clk), .Q(\mem[8][17] ) );
  DFFX1 \mem_reg[8][16]  ( .D(n386), .CLK(clk), .Q(\mem[8][16] ) );
  DFFX1 \mem_reg[8][15]  ( .D(n385), .CLK(clk), .Q(\mem[8][15] ) );
  DFFX1 \mem_reg[8][14]  ( .D(n384), .CLK(clk), .Q(\mem[8][14] ) );
  DFFX1 \mem_reg[8][13]  ( .D(n383), .CLK(clk), .Q(\mem[8][13] ) );
  DFFX1 \mem_reg[8][12]  ( .D(n382), .CLK(clk), .Q(\mem[8][12] ) );
  DFFX1 \mem_reg[8][11]  ( .D(n381), .CLK(clk), .Q(\mem[8][11] ) );
  DFFX1 \mem_reg[8][10]  ( .D(n380), .CLK(clk), .Q(\mem[8][10] ) );
  DFFX1 \mem_reg[8][9]  ( .D(n379), .CLK(clk), .Q(\mem[8][9] ) );
  DFFX1 \mem_reg[8][8]  ( .D(n378), .CLK(clk), .Q(\mem[8][8] ) );
  DFFX1 \mem_reg[8][7]  ( .D(n377), .CLK(clk), .Q(\mem[8][7] ) );
  DFFX1 \mem_reg[8][6]  ( .D(n376), .CLK(clk), .Q(\mem[8][6] ) );
  DFFX1 \mem_reg[8][5]  ( .D(n375), .CLK(clk), .Q(\mem[8][5] ) );
  DFFX1 \mem_reg[8][4]  ( .D(n374), .CLK(clk), .Q(\mem[8][4] ) );
  DFFX1 \mem_reg[8][3]  ( .D(n373), .CLK(clk), .Q(\mem[8][3] ) );
  DFFX1 \mem_reg[8][2]  ( .D(n372), .CLK(clk), .Q(\mem[8][2] ) );
  DFFX1 \mem_reg[8][1]  ( .D(n371), .CLK(clk), .Q(\mem[8][1] ) );
  DFFX1 \mem_reg[8][0]  ( .D(n370), .CLK(clk), .Q(\mem[8][0] ) );
  DFFX1 \mem_reg[7][31]  ( .D(n369), .CLK(clk), .Q(\mem[7][31] ) );
  DFFX1 \mem_reg[7][30]  ( .D(n368), .CLK(clk), .Q(\mem[7][30] ) );
  DFFX1 \mem_reg[7][29]  ( .D(n367), .CLK(clk), .Q(\mem[7][29] ) );
  DFFX1 \mem_reg[7][28]  ( .D(n366), .CLK(clk), .Q(\mem[7][28] ) );
  DFFX1 \mem_reg[7][27]  ( .D(n365), .CLK(clk), .Q(\mem[7][27] ) );
  DFFX1 \mem_reg[7][26]  ( .D(n364), .CLK(clk), .Q(\mem[7][26] ) );
  DFFX1 \mem_reg[7][25]  ( .D(n363), .CLK(clk), .Q(\mem[7][25] ) );
  DFFX1 \mem_reg[7][24]  ( .D(n362), .CLK(clk), .Q(\mem[7][24] ) );
  DFFX1 \mem_reg[7][23]  ( .D(n361), .CLK(clk), .Q(\mem[7][23] ) );
  DFFX1 \mem_reg[7][22]  ( .D(n360), .CLK(clk), .Q(\mem[7][22] ) );
  DFFX1 \mem_reg[7][21]  ( .D(n359), .CLK(clk), .Q(\mem[7][21] ) );
  DFFX1 \mem_reg[7][20]  ( .D(n358), .CLK(clk), .Q(\mem[7][20] ) );
  DFFX1 \mem_reg[7][19]  ( .D(n357), .CLK(clk), .Q(\mem[7][19] ) );
  DFFX1 \mem_reg[7][18]  ( .D(n356), .CLK(clk), .Q(\mem[7][18] ) );
  DFFX1 \mem_reg[7][17]  ( .D(n355), .CLK(clk), .Q(\mem[7][17] ) );
  DFFX1 \mem_reg[7][16]  ( .D(n354), .CLK(clk), .Q(\mem[7][16] ) );
  DFFX1 \mem_reg[7][15]  ( .D(n353), .CLK(clk), .Q(\mem[7][15] ) );
  DFFX1 \mem_reg[7][14]  ( .D(n352), .CLK(clk), .Q(\mem[7][14] ) );
  DFFX1 \mem_reg[7][13]  ( .D(n351), .CLK(clk), .Q(\mem[7][13] ) );
  DFFX1 \mem_reg[7][12]  ( .D(n350), .CLK(clk), .Q(\mem[7][12] ) );
  DFFX1 \mem_reg[7][11]  ( .D(n349), .CLK(clk), .Q(\mem[7][11] ) );
  DFFX1 \mem_reg[7][10]  ( .D(n348), .CLK(clk), .Q(\mem[7][10] ) );
  DFFX1 \mem_reg[7][9]  ( .D(n347), .CLK(clk), .Q(\mem[7][9] ) );
  DFFX1 \mem_reg[7][8]  ( .D(n346), .CLK(clk), .Q(\mem[7][8] ) );
  DFFX1 \mem_reg[7][7]  ( .D(n345), .CLK(clk), .Q(\mem[7][7] ) );
  DFFX1 \mem_reg[7][6]  ( .D(n344), .CLK(clk), .Q(\mem[7][6] ) );
  DFFX1 \mem_reg[7][5]  ( .D(n343), .CLK(clk), .Q(\mem[7][5] ) );
  DFFX1 \mem_reg[7][4]  ( .D(n342), .CLK(clk), .Q(\mem[7][4] ) );
  DFFX1 \mem_reg[7][3]  ( .D(n341), .CLK(clk), .Q(\mem[7][3] ) );
  DFFX1 \mem_reg[7][2]  ( .D(n340), .CLK(clk), .Q(\mem[7][2] ) );
  DFFX1 \mem_reg[7][1]  ( .D(n339), .CLK(clk), .Q(\mem[7][1] ) );
  DFFX1 \mem_reg[7][0]  ( .D(n338), .CLK(clk), .Q(\mem[7][0] ) );
  DFFX1 \mem_reg[6][31]  ( .D(n337), .CLK(clk), .Q(\mem[6][31] ) );
  DFFX1 \mem_reg[6][30]  ( .D(n336), .CLK(clk), .Q(\mem[6][30] ) );
  DFFX1 \mem_reg[6][29]  ( .D(n335), .CLK(clk), .Q(\mem[6][29] ) );
  DFFX1 \mem_reg[6][28]  ( .D(n334), .CLK(clk), .Q(\mem[6][28] ) );
  DFFX1 \mem_reg[6][27]  ( .D(n333), .CLK(clk), .Q(\mem[6][27] ) );
  DFFX1 \mem_reg[6][26]  ( .D(n332), .CLK(clk), .Q(\mem[6][26] ) );
  DFFX1 \mem_reg[6][25]  ( .D(n331), .CLK(clk), .Q(\mem[6][25] ) );
  DFFX1 \mem_reg[6][24]  ( .D(n330), .CLK(clk), .Q(\mem[6][24] ) );
  DFFX1 \mem_reg[6][23]  ( .D(n329), .CLK(clk), .Q(\mem[6][23] ) );
  DFFX1 \mem_reg[6][22]  ( .D(n328), .CLK(clk), .Q(\mem[6][22] ) );
  DFFX1 \mem_reg[6][21]  ( .D(n327), .CLK(clk), .Q(\mem[6][21] ) );
  DFFX1 \mem_reg[6][20]  ( .D(n326), .CLK(clk), .Q(\mem[6][20] ) );
  DFFX1 \mem_reg[6][19]  ( .D(n325), .CLK(clk), .Q(\mem[6][19] ) );
  DFFX1 \mem_reg[6][18]  ( .D(n324), .CLK(clk), .Q(\mem[6][18] ) );
  DFFX1 \mem_reg[6][17]  ( .D(n323), .CLK(clk), .Q(\mem[6][17] ) );
  DFFX1 \mem_reg[6][16]  ( .D(n322), .CLK(clk), .Q(\mem[6][16] ) );
  DFFX1 \mem_reg[6][15]  ( .D(n321), .CLK(clk), .Q(\mem[6][15] ) );
  DFFX1 \mem_reg[6][14]  ( .D(n320), .CLK(clk), .Q(\mem[6][14] ) );
  DFFX1 \mem_reg[6][13]  ( .D(n319), .CLK(clk), .Q(\mem[6][13] ) );
  DFFX1 \mem_reg[6][12]  ( .D(n318), .CLK(clk), .Q(\mem[6][12] ) );
  DFFX1 \mem_reg[6][11]  ( .D(n317), .CLK(clk), .Q(\mem[6][11] ) );
  DFFX1 \mem_reg[6][10]  ( .D(n316), .CLK(clk), .Q(\mem[6][10] ) );
  DFFX1 \mem_reg[6][9]  ( .D(n315), .CLK(clk), .Q(\mem[6][9] ) );
  DFFX1 \mem_reg[6][8]  ( .D(n314), .CLK(clk), .Q(\mem[6][8] ) );
  DFFX1 \mem_reg[6][7]  ( .D(n313), .CLK(clk), .Q(\mem[6][7] ) );
  DFFX1 \mem_reg[6][6]  ( .D(n312), .CLK(clk), .Q(\mem[6][6] ) );
  DFFX1 \mem_reg[6][5]  ( .D(n311), .CLK(clk), .Q(\mem[6][5] ) );
  DFFX1 \mem_reg[6][4]  ( .D(n310), .CLK(clk), .Q(\mem[6][4] ) );
  DFFX1 \mem_reg[6][3]  ( .D(n309), .CLK(clk), .Q(\mem[6][3] ) );
  DFFX1 \mem_reg[6][2]  ( .D(n308), .CLK(clk), .Q(\mem[6][2] ) );
  DFFX1 \mem_reg[6][1]  ( .D(n307), .CLK(clk), .Q(\mem[6][1] ) );
  DFFX1 \mem_reg[6][0]  ( .D(n306), .CLK(clk), .Q(\mem[6][0] ) );
  DFFX1 \mem_reg[5][31]  ( .D(n305), .CLK(clk), .Q(\mem[5][31] ) );
  DFFX1 \mem_reg[5][30]  ( .D(n304), .CLK(clk), .Q(\mem[5][30] ) );
  DFFX1 \mem_reg[5][29]  ( .D(n303), .CLK(clk), .Q(\mem[5][29] ) );
  DFFX1 \mem_reg[5][28]  ( .D(n302), .CLK(clk), .Q(\mem[5][28] ) );
  DFFX1 \mem_reg[5][27]  ( .D(n301), .CLK(clk), .Q(\mem[5][27] ) );
  DFFX1 \mem_reg[5][26]  ( .D(n300), .CLK(clk), .Q(\mem[5][26] ) );
  DFFX1 \mem_reg[5][25]  ( .D(n299), .CLK(clk), .Q(\mem[5][25] ) );
  DFFX1 \mem_reg[5][24]  ( .D(n298), .CLK(clk), .Q(\mem[5][24] ) );
  DFFX1 \mem_reg[5][23]  ( .D(n297), .CLK(clk), .Q(\mem[5][23] ) );
  DFFX1 \mem_reg[5][22]  ( .D(n296), .CLK(clk), .Q(\mem[5][22] ) );
  DFFX1 \mem_reg[5][21]  ( .D(n295), .CLK(clk), .Q(\mem[5][21] ) );
  DFFX1 \mem_reg[5][20]  ( .D(n294), .CLK(clk), .Q(\mem[5][20] ) );
  DFFX1 \mem_reg[5][19]  ( .D(n293), .CLK(clk), .Q(\mem[5][19] ) );
  DFFX1 \mem_reg[5][18]  ( .D(n292), .CLK(clk), .Q(\mem[5][18] ) );
  DFFX1 \mem_reg[5][17]  ( .D(n291), .CLK(clk), .Q(\mem[5][17] ) );
  DFFX1 \mem_reg[5][16]  ( .D(n290), .CLK(clk), .Q(\mem[5][16] ) );
  DFFX1 \mem_reg[5][15]  ( .D(n289), .CLK(clk), .Q(\mem[5][15] ) );
  DFFX1 \mem_reg[5][14]  ( .D(n288), .CLK(clk), .Q(\mem[5][14] ) );
  DFFX1 \mem_reg[5][13]  ( .D(n287), .CLK(clk), .Q(\mem[5][13] ) );
  DFFX1 \mem_reg[5][12]  ( .D(n286), .CLK(clk), .Q(\mem[5][12] ) );
  DFFX1 \mem_reg[5][11]  ( .D(n285), .CLK(clk), .Q(\mem[5][11] ) );
  DFFX1 \mem_reg[5][10]  ( .D(n284), .CLK(clk), .Q(\mem[5][10] ) );
  DFFX1 \mem_reg[5][9]  ( .D(n283), .CLK(clk), .Q(\mem[5][9] ) );
  DFFX1 \mem_reg[5][8]  ( .D(n282), .CLK(clk), .Q(\mem[5][8] ) );
  DFFX1 \mem_reg[5][7]  ( .D(n281), .CLK(clk), .Q(\mem[5][7] ) );
  DFFX1 \mem_reg[5][6]  ( .D(n280), .CLK(clk), .Q(\mem[5][6] ) );
  DFFX1 \mem_reg[5][5]  ( .D(n279), .CLK(clk), .Q(\mem[5][5] ) );
  DFFX1 \mem_reg[5][4]  ( .D(n278), .CLK(clk), .Q(\mem[5][4] ) );
  DFFX1 \mem_reg[5][3]  ( .D(n277), .CLK(clk), .Q(\mem[5][3] ) );
  DFFX1 \mem_reg[5][2]  ( .D(n276), .CLK(clk), .Q(\mem[5][2] ) );
  DFFX1 \mem_reg[5][1]  ( .D(n275), .CLK(clk), .Q(\mem[5][1] ) );
  DFFX1 \mem_reg[5][0]  ( .D(n274), .CLK(clk), .Q(\mem[5][0] ) );
  DFFX1 \mem_reg[4][31]  ( .D(n273), .CLK(clk), .Q(\mem[4][31] ) );
  DFFX1 \mem_reg[4][30]  ( .D(n272), .CLK(clk), .Q(\mem[4][30] ) );
  DFFX1 \mem_reg[4][29]  ( .D(n271), .CLK(clk), .Q(\mem[4][29] ) );
  DFFX1 \mem_reg[4][28]  ( .D(n270), .CLK(clk), .Q(\mem[4][28] ) );
  DFFX1 \mem_reg[4][27]  ( .D(n269), .CLK(clk), .Q(\mem[4][27] ) );
  DFFX1 \mem_reg[4][26]  ( .D(n268), .CLK(clk), .Q(\mem[4][26] ) );
  DFFX1 \mem_reg[4][25]  ( .D(n267), .CLK(clk), .Q(\mem[4][25] ) );
  DFFX1 \mem_reg[4][24]  ( .D(n266), .CLK(clk), .Q(\mem[4][24] ) );
  DFFX1 \mem_reg[4][23]  ( .D(n265), .CLK(clk), .Q(\mem[4][23] ) );
  DFFX1 \mem_reg[4][22]  ( .D(n264), .CLK(clk), .Q(\mem[4][22] ) );
  DFFX1 \mem_reg[4][21]  ( .D(n263), .CLK(clk), .Q(\mem[4][21] ) );
  DFFX1 \mem_reg[4][20]  ( .D(n262), .CLK(clk), .Q(\mem[4][20] ) );
  DFFX1 \mem_reg[4][19]  ( .D(n261), .CLK(clk), .Q(\mem[4][19] ) );
  DFFX1 \mem_reg[4][18]  ( .D(n260), .CLK(clk), .Q(\mem[4][18] ) );
  DFFX1 \mem_reg[4][17]  ( .D(n259), .CLK(clk), .Q(\mem[4][17] ) );
  DFFX1 \mem_reg[4][16]  ( .D(n258), .CLK(clk), .Q(\mem[4][16] ) );
  DFFX1 \mem_reg[4][15]  ( .D(n257), .CLK(clk), .Q(\mem[4][15] ) );
  DFFX1 \mem_reg[4][14]  ( .D(n256), .CLK(clk), .Q(\mem[4][14] ) );
  DFFX1 \mem_reg[4][13]  ( .D(n255), .CLK(clk), .Q(\mem[4][13] ) );
  DFFX1 \mem_reg[4][12]  ( .D(n254), .CLK(clk), .Q(\mem[4][12] ) );
  DFFX1 \mem_reg[4][11]  ( .D(n253), .CLK(clk), .Q(\mem[4][11] ) );
  DFFX1 \mem_reg[4][10]  ( .D(n252), .CLK(clk), .Q(\mem[4][10] ) );
  DFFX1 \mem_reg[4][9]  ( .D(n251), .CLK(clk), .Q(\mem[4][9] ) );
  DFFX1 \mem_reg[4][8]  ( .D(n250), .CLK(clk), .Q(\mem[4][8] ) );
  DFFX1 \mem_reg[4][7]  ( .D(n249), .CLK(clk), .Q(\mem[4][7] ) );
  DFFX1 \mem_reg[4][6]  ( .D(n248), .CLK(clk), .Q(\mem[4][6] ) );
  DFFX1 \mem_reg[4][5]  ( .D(n247), .CLK(clk), .Q(\mem[4][5] ) );
  DFFX1 \mem_reg[4][4]  ( .D(n246), .CLK(clk), .Q(\mem[4][4] ) );
  DFFX1 \mem_reg[4][3]  ( .D(n245), .CLK(clk), .Q(\mem[4][3] ) );
  DFFX1 \mem_reg[4][2]  ( .D(n244), .CLK(clk), .Q(\mem[4][2] ) );
  DFFX1 \mem_reg[4][1]  ( .D(n243), .CLK(clk), .Q(\mem[4][1] ) );
  DFFX1 \mem_reg[4][0]  ( .D(n242), .CLK(clk), .Q(\mem[4][0] ) );
  DFFX1 \mem_reg[3][31]  ( .D(n241), .CLK(clk), .Q(\mem[3][31] ) );
  DFFX1 \mem_reg[3][30]  ( .D(n240), .CLK(clk), .Q(\mem[3][30] ) );
  DFFX1 \mem_reg[3][29]  ( .D(n239), .CLK(clk), .Q(\mem[3][29] ) );
  DFFX1 \mem_reg[3][28]  ( .D(n238), .CLK(clk), .Q(\mem[3][28] ) );
  DFFX1 \mem_reg[3][27]  ( .D(n237), .CLK(clk), .Q(\mem[3][27] ) );
  DFFX1 \mem_reg[3][26]  ( .D(n236), .CLK(clk), .Q(\mem[3][26] ) );
  DFFX1 \mem_reg[3][25]  ( .D(n235), .CLK(clk), .Q(\mem[3][25] ) );
  DFFX1 \mem_reg[3][24]  ( .D(n234), .CLK(clk), .Q(\mem[3][24] ) );
  DFFX1 \mem_reg[3][23]  ( .D(n233), .CLK(clk), .Q(\mem[3][23] ) );
  DFFX1 \mem_reg[3][22]  ( .D(n232), .CLK(clk), .Q(\mem[3][22] ) );
  DFFX1 \mem_reg[3][21]  ( .D(n231), .CLK(clk), .Q(\mem[3][21] ) );
  DFFX1 \mem_reg[3][20]  ( .D(n230), .CLK(clk), .Q(\mem[3][20] ) );
  DFFX1 \mem_reg[3][19]  ( .D(n229), .CLK(clk), .Q(\mem[3][19] ) );
  DFFX1 \mem_reg[3][18]  ( .D(n228), .CLK(clk), .Q(\mem[3][18] ) );
  DFFX1 \mem_reg[3][17]  ( .D(n227), .CLK(clk), .Q(\mem[3][17] ) );
  DFFX1 \mem_reg[3][16]  ( .D(n226), .CLK(clk), .Q(\mem[3][16] ) );
  DFFX1 \mem_reg[3][15]  ( .D(n225), .CLK(clk), .Q(\mem[3][15] ) );
  DFFX1 \mem_reg[3][14]  ( .D(n224), .CLK(clk), .Q(\mem[3][14] ) );
  DFFX1 \mem_reg[3][13]  ( .D(n223), .CLK(clk), .Q(\mem[3][13] ) );
  DFFX1 \mem_reg[3][12]  ( .D(n222), .CLK(clk), .Q(\mem[3][12] ) );
  DFFX1 \mem_reg[3][11]  ( .D(n221), .CLK(clk), .Q(\mem[3][11] ) );
  DFFX1 \mem_reg[3][10]  ( .D(n220), .CLK(clk), .Q(\mem[3][10] ) );
  DFFX1 \mem_reg[3][9]  ( .D(n219), .CLK(clk), .Q(\mem[3][9] ) );
  DFFX1 \mem_reg[3][8]  ( .D(n218), .CLK(clk), .Q(\mem[3][8] ) );
  DFFX1 \mem_reg[3][7]  ( .D(n217), .CLK(clk), .Q(\mem[3][7] ) );
  DFFX1 \mem_reg[3][6]  ( .D(n216), .CLK(clk), .Q(\mem[3][6] ) );
  DFFX1 \mem_reg[3][5]  ( .D(n215), .CLK(clk), .Q(\mem[3][5] ) );
  DFFX1 \mem_reg[3][4]  ( .D(n214), .CLK(clk), .Q(\mem[3][4] ) );
  DFFX1 \mem_reg[3][3]  ( .D(n213), .CLK(clk), .Q(\mem[3][3] ) );
  DFFX1 \mem_reg[3][2]  ( .D(n212), .CLK(clk), .Q(\mem[3][2] ) );
  DFFX1 \mem_reg[3][1]  ( .D(n211), .CLK(clk), .Q(\mem[3][1] ) );
  DFFX1 \mem_reg[3][0]  ( .D(n210), .CLK(clk), .Q(\mem[3][0] ) );
  DFFX1 \mem_reg[2][31]  ( .D(n209), .CLK(clk), .Q(\mem[2][31] ) );
  DFFX1 \mem_reg[2][30]  ( .D(n208), .CLK(clk), .Q(\mem[2][30] ) );
  DFFX1 \mem_reg[2][29]  ( .D(n207), .CLK(clk), .Q(\mem[2][29] ) );
  DFFX1 \mem_reg[2][28]  ( .D(n206), .CLK(clk), .Q(\mem[2][28] ) );
  DFFX1 \mem_reg[2][27]  ( .D(n205), .CLK(clk), .Q(\mem[2][27] ) );
  DFFX1 \mem_reg[2][26]  ( .D(n204), .CLK(clk), .Q(\mem[2][26] ) );
  DFFX1 \mem_reg[2][25]  ( .D(n203), .CLK(clk), .Q(\mem[2][25] ) );
  DFFX1 \mem_reg[2][24]  ( .D(n202), .CLK(clk), .Q(\mem[2][24] ) );
  DFFX1 \mem_reg[2][23]  ( .D(n201), .CLK(clk), .Q(\mem[2][23] ) );
  DFFX1 \mem_reg[2][22]  ( .D(n200), .CLK(clk), .Q(\mem[2][22] ) );
  DFFX1 \mem_reg[2][21]  ( .D(n199), .CLK(clk), .Q(\mem[2][21] ) );
  DFFX1 \mem_reg[2][20]  ( .D(n198), .CLK(clk), .Q(\mem[2][20] ) );
  DFFX1 \mem_reg[2][19]  ( .D(n197), .CLK(clk), .Q(\mem[2][19] ) );
  DFFX1 \mem_reg[2][18]  ( .D(n196), .CLK(clk), .Q(\mem[2][18] ) );
  DFFX1 \mem_reg[2][17]  ( .D(n195), .CLK(clk), .Q(\mem[2][17] ) );
  DFFX1 \mem_reg[2][16]  ( .D(n194), .CLK(clk), .Q(\mem[2][16] ) );
  DFFX1 \mem_reg[2][15]  ( .D(n193), .CLK(clk), .Q(\mem[2][15] ) );
  DFFX1 \mem_reg[2][14]  ( .D(n192), .CLK(clk), .Q(\mem[2][14] ) );
  DFFX1 \mem_reg[2][13]  ( .D(n191), .CLK(clk), .Q(\mem[2][13] ) );
  DFFX1 \mem_reg[2][12]  ( .D(n190), .CLK(clk), .Q(\mem[2][12] ) );
  DFFX1 \mem_reg[2][11]  ( .D(n189), .CLK(clk), .Q(\mem[2][11] ) );
  DFFX1 \mem_reg[2][10]  ( .D(n188), .CLK(clk), .Q(\mem[2][10] ) );
  DFFX1 \mem_reg[2][9]  ( .D(n187), .CLK(clk), .Q(\mem[2][9] ) );
  DFFX1 \mem_reg[2][8]  ( .D(n186), .CLK(clk), .Q(\mem[2][8] ) );
  DFFX1 \mem_reg[2][7]  ( .D(n185), .CLK(clk), .Q(\mem[2][7] ) );
  DFFX1 \mem_reg[2][6]  ( .D(n184), .CLK(clk), .Q(\mem[2][6] ) );
  DFFX1 \mem_reg[2][5]  ( .D(n183), .CLK(clk), .Q(\mem[2][5] ) );
  DFFX1 \mem_reg[2][4]  ( .D(n182), .CLK(clk), .Q(\mem[2][4] ) );
  DFFX1 \mem_reg[2][3]  ( .D(n181), .CLK(clk), .Q(\mem[2][3] ) );
  DFFX1 \mem_reg[2][2]  ( .D(n180), .CLK(clk), .Q(\mem[2][2] ) );
  DFFX1 \mem_reg[2][1]  ( .D(n179), .CLK(clk), .Q(\mem[2][1] ) );
  DFFX1 \mem_reg[2][0]  ( .D(n178), .CLK(clk), .Q(\mem[2][0] ) );
  DFFX1 \mem_reg[1][31]  ( .D(n177), .CLK(clk), .Q(\mem[1][31] ) );
  DFFX1 \mem_reg[1][30]  ( .D(n176), .CLK(clk), .Q(\mem[1][30] ) );
  DFFX1 \mem_reg[1][29]  ( .D(n175), .CLK(clk), .Q(\mem[1][29] ) );
  DFFX1 \mem_reg[1][28]  ( .D(n174), .CLK(clk), .Q(\mem[1][28] ) );
  DFFX1 \mem_reg[1][27]  ( .D(n173), .CLK(clk), .Q(\mem[1][27] ) );
  DFFX1 \mem_reg[1][26]  ( .D(n172), .CLK(clk), .Q(\mem[1][26] ) );
  DFFX1 \mem_reg[1][25]  ( .D(n171), .CLK(clk), .Q(\mem[1][25] ) );
  DFFX1 \mem_reg[1][24]  ( .D(n170), .CLK(clk), .Q(\mem[1][24] ) );
  DFFX1 \mem_reg[1][23]  ( .D(n169), .CLK(clk), .Q(\mem[1][23] ) );
  DFFX1 \mem_reg[1][22]  ( .D(n168), .CLK(clk), .Q(\mem[1][22] ) );
  DFFX1 \mem_reg[1][21]  ( .D(n167), .CLK(clk), .Q(\mem[1][21] ) );
  DFFX1 \mem_reg[1][20]  ( .D(n166), .CLK(clk), .Q(\mem[1][20] ) );
  DFFX1 \mem_reg[1][19]  ( .D(n165), .CLK(clk), .Q(\mem[1][19] ) );
  DFFX1 \mem_reg[1][18]  ( .D(n164), .CLK(clk), .Q(\mem[1][18] ) );
  DFFX1 \mem_reg[1][17]  ( .D(n163), .CLK(clk), .Q(\mem[1][17] ) );
  DFFX1 \mem_reg[1][16]  ( .D(n162), .CLK(clk), .Q(\mem[1][16] ) );
  DFFX1 \mem_reg[1][15]  ( .D(n161), .CLK(clk), .Q(\mem[1][15] ) );
  DFFX1 \mem_reg[1][14]  ( .D(n160), .CLK(clk), .Q(\mem[1][14] ) );
  DFFX1 \mem_reg[1][13]  ( .D(n159), .CLK(clk), .Q(\mem[1][13] ) );
  DFFX1 \mem_reg[1][12]  ( .D(n158), .CLK(clk), .Q(\mem[1][12] ) );
  DFFX1 \mem_reg[1][11]  ( .D(n157), .CLK(clk), .Q(\mem[1][11] ) );
  DFFX1 \mem_reg[1][10]  ( .D(n156), .CLK(clk), .Q(\mem[1][10] ) );
  DFFX1 \mem_reg[1][9]  ( .D(n155), .CLK(clk), .Q(\mem[1][9] ) );
  DFFX1 \mem_reg[1][8]  ( .D(n154), .CLK(clk), .Q(\mem[1][8] ) );
  DFFX1 \mem_reg[1][7]  ( .D(n153), .CLK(clk), .Q(\mem[1][7] ) );
  DFFX1 \mem_reg[1][6]  ( .D(n152), .CLK(clk), .Q(\mem[1][6] ) );
  DFFX1 \mem_reg[1][5]  ( .D(n151), .CLK(clk), .Q(\mem[1][5] ) );
  DFFX1 \mem_reg[1][4]  ( .D(n150), .CLK(clk), .Q(\mem[1][4] ) );
  DFFX1 \mem_reg[1][3]  ( .D(n149), .CLK(clk), .Q(\mem[1][3] ) );
  DFFX1 \mem_reg[1][2]  ( .D(n148), .CLK(clk), .Q(\mem[1][2] ) );
  DFFX1 \mem_reg[1][1]  ( .D(n147), .CLK(clk), .Q(\mem[1][1] ) );
  DFFX1 \mem_reg[1][0]  ( .D(n146), .CLK(clk), .Q(\mem[1][0] ) );
  DFFX1 \mem_reg[0][31]  ( .D(n145), .CLK(clk), .Q(\mem[0][31] ) );
  DFFX1 \mem_reg[0][30]  ( .D(n144), .CLK(clk), .Q(\mem[0][30] ) );
  DFFX1 \mem_reg[0][29]  ( .D(n143), .CLK(clk), .Q(\mem[0][29] ) );
  DFFX1 \mem_reg[0][28]  ( .D(n142), .CLK(clk), .Q(\mem[0][28] ) );
  DFFX1 \mem_reg[0][27]  ( .D(n141), .CLK(clk), .Q(\mem[0][27] ) );
  DFFX1 \mem_reg[0][26]  ( .D(n140), .CLK(clk), .Q(\mem[0][26] ) );
  DFFX1 \mem_reg[0][25]  ( .D(n139), .CLK(clk), .Q(\mem[0][25] ) );
  DFFX1 \mem_reg[0][24]  ( .D(n138), .CLK(clk), .Q(\mem[0][24] ) );
  DFFX1 \mem_reg[0][23]  ( .D(n137), .CLK(clk), .Q(\mem[0][23] ) );
  DFFX1 \mem_reg[0][22]  ( .D(n136), .CLK(clk), .Q(\mem[0][22] ) );
  DFFX1 \mem_reg[0][21]  ( .D(n135), .CLK(clk), .Q(\mem[0][21] ) );
  DFFX1 \mem_reg[0][20]  ( .D(n134), .CLK(clk), .Q(\mem[0][20] ) );
  DFFX1 \mem_reg[0][19]  ( .D(n133), .CLK(clk), .Q(\mem[0][19] ) );
  DFFX1 \mem_reg[0][18]  ( .D(n132), .CLK(clk), .Q(\mem[0][18] ) );
  DFFX1 \mem_reg[0][17]  ( .D(n131), .CLK(clk), .Q(\mem[0][17] ) );
  DFFX1 \mem_reg[0][16]  ( .D(n130), .CLK(clk), .Q(\mem[0][16] ) );
  DFFX1 \mem_reg[0][15]  ( .D(n129), .CLK(clk), .Q(\mem[0][15] ) );
  DFFX1 \mem_reg[0][14]  ( .D(n128), .CLK(clk), .Q(\mem[0][14] ) );
  DFFX1 \mem_reg[0][13]  ( .D(n127), .CLK(clk), .Q(\mem[0][13] ) );
  DFFX1 \mem_reg[0][12]  ( .D(n126), .CLK(clk), .Q(\mem[0][12] ) );
  DFFX1 \mem_reg[0][11]  ( .D(n125), .CLK(clk), .Q(\mem[0][11] ) );
  DFFX1 \mem_reg[0][10]  ( .D(n124), .CLK(clk), .Q(\mem[0][10] ) );
  DFFX1 \mem_reg[0][9]  ( .D(n123), .CLK(clk), .Q(\mem[0][9] ) );
  DFFX1 \mem_reg[0][8]  ( .D(n122), .CLK(clk), .Q(\mem[0][8] ) );
  DFFX1 \mem_reg[0][7]  ( .D(n121), .CLK(clk), .Q(\mem[0][7] ) );
  DFFX1 \mem_reg[0][6]  ( .D(n120), .CLK(clk), .Q(\mem[0][6] ) );
  DFFX1 \mem_reg[0][5]  ( .D(n119), .CLK(clk), .Q(\mem[0][5] ) );
  DFFX1 \mem_reg[0][4]  ( .D(n118), .CLK(clk), .Q(\mem[0][4] ) );
  DFFX1 \mem_reg[0][3]  ( .D(n117), .CLK(clk), .Q(\mem[0][3] ) );
  DFFX1 \mem_reg[0][2]  ( .D(n116), .CLK(clk), .Q(\mem[0][2] ) );
  DFFX1 \mem_reg[0][1]  ( .D(n115), .CLK(clk), .Q(\mem[0][1] ) );
  DFFX1 \mem_reg[0][0]  ( .D(n114), .CLK(clk), .Q(\mem[0][0] ) );
  AO22X1 U40 ( .IN1(n1875), .IN2(n1842), .IN3(\mem[26][13] ), .IN4(n1995), .Q(
        n959) );
  AO22X1 U41 ( .IN1(n1873), .IN2(n1841), .IN3(\mem[26][14] ), .IN4(n1995), .Q(
        n960) );
  AO22X1 U42 ( .IN1(n1871), .IN2(n39), .IN3(\mem[26][15] ), .IN4(n1995), .Q(
        n961) );
  AO22X1 U43 ( .IN1(n1869), .IN2(n1842), .IN3(\mem[26][16] ), .IN4(n1995), .Q(
        n962) );
  AO22X1 U44 ( .IN1(n1867), .IN2(n1841), .IN3(\mem[26][17] ), .IN4(n1995), .Q(
        n963) );
  AO22X1 U45 ( .IN1(n1865), .IN2(n39), .IN3(\mem[26][18] ), .IN4(n1995), .Q(
        n964) );
  AO22X1 U46 ( .IN1(n1863), .IN2(n1842), .IN3(\mem[26][19] ), .IN4(n1995), .Q(
        n965) );
  AO22X1 U47 ( .IN1(n1861), .IN2(n1841), .IN3(\mem[26][20] ), .IN4(n1995), .Q(
        n966) );
  AO22X1 U48 ( .IN1(n1859), .IN2(n39), .IN3(\mem[26][21] ), .IN4(n1995), .Q(
        n967) );
  AO22X1 U49 ( .IN1(n1857), .IN2(n1842), .IN3(\mem[26][22] ), .IN4(n1995), .Q(
        n968) );
  AO22X1 U50 ( .IN1(n1855), .IN2(n1841), .IN3(\mem[26][23] ), .IN4(n1995), .Q(
        n969) );
  AO22X1 U51 ( .IN1(n1854), .IN2(n39), .IN3(\mem[26][24] ), .IN4(n1995), .Q(
        n970) );
  AO22X1 U52 ( .IN1(n1853), .IN2(n1842), .IN3(\mem[26][25] ), .IN4(n1996), .Q(
        n971) );
  AO22X1 U53 ( .IN1(n1852), .IN2(n1841), .IN3(\mem[26][26] ), .IN4(n1996), .Q(
        n972) );
  AO22X1 U54 ( .IN1(n1851), .IN2(n39), .IN3(\mem[26][27] ), .IN4(n1996), .Q(
        n973) );
  AO22X1 U55 ( .IN1(n1850), .IN2(n1842), .IN3(\mem[26][28] ), .IN4(n1996), .Q(
        n974) );
  AO22X1 U56 ( .IN1(n1849), .IN2(n1841), .IN3(\mem[26][29] ), .IN4(n1996), .Q(
        n975) );
  AO22X1 U57 ( .IN1(n1848), .IN2(n39), .IN3(\mem[26][30] ), .IN4(n1996), .Q(
        n976) );
  AO22X1 U58 ( .IN1(n1845), .IN2(n1842), .IN3(\mem[26][31] ), .IN4(n1996), .Q(
        n977) );
  AO22X1 U59 ( .IN1(n1844), .IN2(n1934), .IN3(\mem[27][0] ), .IN4(n1993), .Q(
        n978) );
  AO22X1 U60 ( .IN1(n1843), .IN2(n1933), .IN3(\mem[27][1] ), .IN4(n1993), .Q(
        n979) );
  AO22X1 U61 ( .IN1(n61), .IN2(n59), .IN3(\mem[27][2] ), .IN4(n1993), .Q(n980)
         );
  AO22X1 U62 ( .IN1(n62), .IN2(n1934), .IN3(\mem[27][3] ), .IN4(n1993), .Q(
        n981) );
  AO22X1 U63 ( .IN1(n63), .IN2(n1933), .IN3(\mem[27][4] ), .IN4(n1993), .Q(
        n982) );
  AO22X1 U64 ( .IN1(n64), .IN2(n59), .IN3(\mem[27][5] ), .IN4(n1993), .Q(n983)
         );
  AO22X1 U65 ( .IN1(n65), .IN2(n1934), .IN3(\mem[27][6] ), .IN4(n1993), .Q(
        n984) );
  AO22X1 U66 ( .IN1(n66), .IN2(n1933), .IN3(\mem[27][7] ), .IN4(n1993), .Q(
        n985) );
  AO22X1 U67 ( .IN1(n67), .IN2(n59), .IN3(\mem[27][8] ), .IN4(n1993), .Q(n986)
         );
  AO22X1 U68 ( .IN1(n68), .IN2(n1934), .IN3(\mem[27][9] ), .IN4(n1993), .Q(
        n987) );
  AO22X1 U69 ( .IN1(n69), .IN2(n1933), .IN3(\mem[27][10] ), .IN4(n1993), .Q(
        n988) );
  AO22X1 U70 ( .IN1(n70), .IN2(n59), .IN3(\mem[27][11] ), .IN4(n1993), .Q(n989) );
  AO22X1 U71 ( .IN1(n71), .IN2(n1934), .IN3(\mem[27][12] ), .IN4(n1994), .Q(
        n990) );
  AO22X1 U72 ( .IN1(n38), .IN2(n1933), .IN3(\mem[27][13] ), .IN4(n1994), .Q(
        n991) );
  AO22X1 U73 ( .IN1(n40), .IN2(n59), .IN3(\mem[27][14] ), .IN4(n1994), .Q(n992) );
  AO22X1 U74 ( .IN1(n41), .IN2(n1934), .IN3(\mem[27][15] ), .IN4(n1994), .Q(
        n993) );
  AO22X1 U75 ( .IN1(n42), .IN2(n1933), .IN3(\mem[27][16] ), .IN4(n1994), .Q(
        n994) );
  AO22X1 U76 ( .IN1(n43), .IN2(n59), .IN3(\mem[27][17] ), .IN4(n1994), .Q(n995) );
  AO22X1 U77 ( .IN1(n44), .IN2(n1934), .IN3(\mem[27][18] ), .IN4(n1994), .Q(
        n996) );
  AO22X1 U78 ( .IN1(n45), .IN2(n1933), .IN3(\mem[27][19] ), .IN4(n1994), .Q(
        n997) );
  AO22X1 U79 ( .IN1(n46), .IN2(n59), .IN3(\mem[27][20] ), .IN4(n1994), .Q(n998) );
  AO22X1 U80 ( .IN1(n47), .IN2(n1934), .IN3(\mem[27][21] ), .IN4(n1994), .Q(
        n999) );
  AO22X1 U81 ( .IN1(n48), .IN2(n1933), .IN3(\mem[27][22] ), .IN4(n1994), .Q(
        n1000) );
  AO22X1 U82 ( .IN1(n49), .IN2(n59), .IN3(\mem[27][23] ), .IN4(n1994), .Q(
        n1001) );
  AO22X1 U83 ( .IN1(n50), .IN2(n1934), .IN3(\mem[27][24] ), .IN4(n1994), .Q(
        n1002) );
  AO22X1 U84 ( .IN1(n51), .IN2(n1933), .IN3(\mem[27][25] ), .IN4(n1994), .Q(
        n1003) );
  AO22X1 U85 ( .IN1(n52), .IN2(n1934), .IN3(\mem[27][26] ), .IN4(n1993), .Q(
        n1004) );
  AO22X1 U86 ( .IN1(n53), .IN2(n1933), .IN3(\mem[27][27] ), .IN4(n1993), .Q(
        n1005) );
  AO22X1 U87 ( .IN1(n54), .IN2(n1934), .IN3(\mem[27][28] ), .IN4(n1994), .Q(
        n1006) );
  AO22X1 U88 ( .IN1(n55), .IN2(n1933), .IN3(\mem[27][29] ), .IN4(n1993), .Q(
        n1007) );
  AO22X1 U89 ( .IN1(n56), .IN2(n1934), .IN3(\mem[27][30] ), .IN4(n1994), .Q(
        n1008) );
  AO22X1 U90 ( .IN1(n57), .IN2(n1933), .IN3(\mem[27][31] ), .IN4(n1993), .Q(
        n1009) );
  AO22X1 U92 ( .IN1(n58), .IN2(n1932), .IN3(\mem[28][0] ), .IN4(n1991), .Q(
        n1010) );
  AO22X1 U93 ( .IN1(n60), .IN2(n1931), .IN3(\mem[28][1] ), .IN4(n1991), .Q(
        n1011) );
  AO22X1 U94 ( .IN1(n61), .IN2(n74), .IN3(\mem[28][2] ), .IN4(n1991), .Q(n1012) );
  AO22X1 U95 ( .IN1(n62), .IN2(n1932), .IN3(\mem[28][3] ), .IN4(n1991), .Q(
        n1013) );
  AO22X1 U96 ( .IN1(n63), .IN2(n1931), .IN3(\mem[28][4] ), .IN4(n1991), .Q(
        n1014) );
  AO22X1 U97 ( .IN1(n64), .IN2(n74), .IN3(\mem[28][5] ), .IN4(n1991), .Q(n1015) );
  AO22X1 U98 ( .IN1(n65), .IN2(n1932), .IN3(\mem[28][6] ), .IN4(n1991), .Q(
        n1016) );
  AO22X1 U99 ( .IN1(n66), .IN2(n1931), .IN3(\mem[28][7] ), .IN4(n1991), .Q(
        n1017) );
  AO22X1 U100 ( .IN1(n67), .IN2(n74), .IN3(\mem[28][8] ), .IN4(n1991), .Q(
        n1018) );
  AO22X1 U101 ( .IN1(n68), .IN2(n1932), .IN3(\mem[28][9] ), .IN4(n1991), .Q(
        n1019) );
  AO22X1 U102 ( .IN1(n69), .IN2(n1931), .IN3(\mem[28][10] ), .IN4(n1991), .Q(
        n1020) );
  AO22X1 U103 ( .IN1(n70), .IN2(n74), .IN3(\mem[28][11] ), .IN4(n1991), .Q(
        n1021) );
  AO22X1 U104 ( .IN1(n71), .IN2(n1932), .IN3(\mem[28][12] ), .IN4(n1992), .Q(
        n1022) );
  AO22X1 U105 ( .IN1(n1876), .IN2(n1931), .IN3(\mem[28][13] ), .IN4(n1992), 
        .Q(n1023) );
  AO22X1 U106 ( .IN1(n1874), .IN2(n74), .IN3(\mem[28][14] ), .IN4(n1992), .Q(
        n1024) );
  AO22X1 U107 ( .IN1(n1872), .IN2(n1932), .IN3(\mem[28][15] ), .IN4(n1992), 
        .Q(n1025) );
  AO22X1 U108 ( .IN1(n1870), .IN2(n1931), .IN3(\mem[28][16] ), .IN4(n1992), 
        .Q(n1026) );
  AO22X1 U109 ( .IN1(n1868), .IN2(n74), .IN3(\mem[28][17] ), .IN4(n1992), .Q(
        n1027) );
  AO22X1 U110 ( .IN1(n1866), .IN2(n1932), .IN3(\mem[28][18] ), .IN4(n1992), 
        .Q(n1028) );
  AO22X1 U111 ( .IN1(n1864), .IN2(n1931), .IN3(\mem[28][19] ), .IN4(n1992), 
        .Q(n1029) );
  AO22X1 U112 ( .IN1(n1862), .IN2(n74), .IN3(\mem[28][20] ), .IN4(n1992), .Q(
        n1030) );
  AO22X1 U113 ( .IN1(n1860), .IN2(n1932), .IN3(\mem[28][21] ), .IN4(n1992), 
        .Q(n1031) );
  AO22X1 U114 ( .IN1(n1858), .IN2(n1931), .IN3(\mem[28][22] ), .IN4(n1992), 
        .Q(n1032) );
  AO22X1 U115 ( .IN1(n1856), .IN2(n74), .IN3(\mem[28][23] ), .IN4(n1992), .Q(
        n1033) );
  AO22X1 U116 ( .IN1(n1854), .IN2(n1932), .IN3(\mem[28][24] ), .IN4(n1992), 
        .Q(n1034) );
  AO22X1 U117 ( .IN1(n1853), .IN2(n1931), .IN3(\mem[28][25] ), .IN4(n1992), 
        .Q(n1035) );
  AO22X1 U118 ( .IN1(n1852), .IN2(n1932), .IN3(\mem[28][26] ), .IN4(n1991), 
        .Q(n1036) );
  AO22X1 U119 ( .IN1(n1851), .IN2(n1931), .IN3(\mem[28][27] ), .IN4(n1992), 
        .Q(n1037) );
  AO22X1 U120 ( .IN1(n1850), .IN2(n1932), .IN3(\mem[28][28] ), .IN4(n1991), 
        .Q(n1038) );
  AO22X1 U121 ( .IN1(n1849), .IN2(n1931), .IN3(\mem[28][29] ), .IN4(n1992), 
        .Q(n1039) );
  AO22X1 U122 ( .IN1(n1848), .IN2(n1932), .IN3(\mem[28][30] ), .IN4(n1991), 
        .Q(n1040) );
  AO22X1 U123 ( .IN1(n1845), .IN2(n1931), .IN3(\mem[28][31] ), .IN4(n1991), 
        .Q(n1041) );
  AO22X1 U125 ( .IN1(n1844), .IN2(n1930), .IN3(\mem[29][0] ), .IN4(n1989), .Q(
        n1042) );
  AO22X1 U126 ( .IN1(n1843), .IN2(n1929), .IN3(\mem[29][1] ), .IN4(n1989), .Q(
        n1043) );
  AO22X1 U127 ( .IN1(n61), .IN2(n76), .IN3(\mem[29][2] ), .IN4(n1989), .Q(
        n1044) );
  AO22X1 U128 ( .IN1(n62), .IN2(n1930), .IN3(\mem[29][3] ), .IN4(n1989), .Q(
        n1045) );
  AO22X1 U129 ( .IN1(n63), .IN2(n1929), .IN3(\mem[29][4] ), .IN4(n1989), .Q(
        n1046) );
  AO22X1 U130 ( .IN1(n64), .IN2(n76), .IN3(\mem[29][5] ), .IN4(n1989), .Q(
        n1047) );
  AO22X1 U131 ( .IN1(n65), .IN2(n1930), .IN3(\mem[29][6] ), .IN4(n1989), .Q(
        n1048) );
  AO22X1 U132 ( .IN1(n66), .IN2(n1929), .IN3(\mem[29][7] ), .IN4(n1989), .Q(
        n1049) );
  AO22X1 U133 ( .IN1(n67), .IN2(n76), .IN3(\mem[29][8] ), .IN4(n1989), .Q(
        n1050) );
  AO22X1 U134 ( .IN1(n68), .IN2(n1930), .IN3(\mem[29][9] ), .IN4(n1989), .Q(
        n1051) );
  AO22X1 U135 ( .IN1(n69), .IN2(n1929), .IN3(\mem[29][10] ), .IN4(n1989), .Q(
        n1052) );
  AO22X1 U136 ( .IN1(n70), .IN2(n76), .IN3(\mem[29][11] ), .IN4(n1989), .Q(
        n1053) );
  AO22X1 U137 ( .IN1(n71), .IN2(n1930), .IN3(\mem[29][12] ), .IN4(n1990), .Q(
        n1054) );
  AO22X1 U138 ( .IN1(n1875), .IN2(n1929), .IN3(\mem[29][13] ), .IN4(n1990), 
        .Q(n1055) );
  AO22X1 U139 ( .IN1(n1873), .IN2(n76), .IN3(\mem[29][14] ), .IN4(n1990), .Q(
        n1056) );
  AO22X1 U140 ( .IN1(n1871), .IN2(n1930), .IN3(\mem[29][15] ), .IN4(n1990), 
        .Q(n1057) );
  AO22X1 U141 ( .IN1(n1869), .IN2(n1929), .IN3(\mem[29][16] ), .IN4(n1990), 
        .Q(n1058) );
  AO22X1 U142 ( .IN1(n1867), .IN2(n76), .IN3(\mem[29][17] ), .IN4(n1990), .Q(
        n1059) );
  AO22X1 U143 ( .IN1(n1865), .IN2(n1930), .IN3(\mem[29][18] ), .IN4(n1990), 
        .Q(n1060) );
  AO22X1 U144 ( .IN1(n1863), .IN2(n1929), .IN3(\mem[29][19] ), .IN4(n1990), 
        .Q(n1061) );
  AO22X1 U145 ( .IN1(n1861), .IN2(n76), .IN3(\mem[29][20] ), .IN4(n1990), .Q(
        n1062) );
  AO22X1 U146 ( .IN1(n1859), .IN2(n1930), .IN3(\mem[29][21] ), .IN4(n1990), 
        .Q(n1063) );
  AO22X1 U147 ( .IN1(n1857), .IN2(n1929), .IN3(\mem[29][22] ), .IN4(n1990), 
        .Q(n1064) );
  AO22X1 U148 ( .IN1(n1855), .IN2(n76), .IN3(\mem[29][23] ), .IN4(n1990), .Q(
        n1065) );
  AO22X1 U149 ( .IN1(n50), .IN2(n1930), .IN3(\mem[29][24] ), .IN4(n1990), .Q(
        n1066) );
  AO22X1 U150 ( .IN1(n51), .IN2(n1929), .IN3(\mem[29][25] ), .IN4(n1990), .Q(
        n1067) );
  AO22X1 U151 ( .IN1(n52), .IN2(n1930), .IN3(\mem[29][26] ), .IN4(n1989), .Q(
        n1068) );
  AO22X1 U152 ( .IN1(n53), .IN2(n1929), .IN3(\mem[29][27] ), .IN4(n1989), .Q(
        n1069) );
  AO22X1 U153 ( .IN1(n54), .IN2(n1930), .IN3(\mem[29][28] ), .IN4(n1990), .Q(
        n1070) );
  AO22X1 U154 ( .IN1(n55), .IN2(n1929), .IN3(\mem[29][29] ), .IN4(n1989), .Q(
        n1071) );
  AO22X1 U155 ( .IN1(n56), .IN2(n1930), .IN3(\mem[29][30] ), .IN4(n1990), .Q(
        n1072) );
  AO22X1 U156 ( .IN1(n57), .IN2(n1929), .IN3(\mem[29][31] ), .IN4(n1989), .Q(
        n1073) );
  AO22X1 U158 ( .IN1(n58), .IN2(n1928), .IN3(\mem[30][0] ), .IN4(n1987), .Q(
        n1074) );
  AO22X1 U159 ( .IN1(n60), .IN2(n1927), .IN3(\mem[30][1] ), .IN4(n1987), .Q(
        n1075) );
  AO22X1 U160 ( .IN1(n61), .IN2(n78), .IN3(\mem[30][2] ), .IN4(n1987), .Q(
        n1076) );
  AO22X1 U161 ( .IN1(n62), .IN2(n1928), .IN3(\mem[30][3] ), .IN4(n1987), .Q(
        n1077) );
  AO22X1 U162 ( .IN1(n63), .IN2(n1927), .IN3(\mem[30][4] ), .IN4(n1987), .Q(
        n1078) );
  AO22X1 U163 ( .IN1(n64), .IN2(n78), .IN3(\mem[30][5] ), .IN4(n1987), .Q(
        n1079) );
  AO22X1 U164 ( .IN1(n65), .IN2(n1928), .IN3(\mem[30][6] ), .IN4(n1987), .Q(
        n1080) );
  AO22X1 U165 ( .IN1(n66), .IN2(n1927), .IN3(\mem[30][7] ), .IN4(n1987), .Q(
        n1081) );
  AO22X1 U166 ( .IN1(n67), .IN2(n78), .IN3(\mem[30][8] ), .IN4(n1987), .Q(
        n1082) );
  AO22X1 U167 ( .IN1(n68), .IN2(n1928), .IN3(\mem[30][9] ), .IN4(n1987), .Q(
        n1083) );
  AO22X1 U168 ( .IN1(n69), .IN2(n1927), .IN3(\mem[30][10] ), .IN4(n1987), .Q(
        n1084) );
  AO22X1 U169 ( .IN1(n70), .IN2(n78), .IN3(\mem[30][11] ), .IN4(n1987), .Q(
        n1085) );
  AO22X1 U170 ( .IN1(n71), .IN2(n1928), .IN3(\mem[30][12] ), .IN4(n1988), .Q(
        n1086) );
  AO22X1 U171 ( .IN1(n38), .IN2(n1927), .IN3(\mem[30][13] ), .IN4(n1988), .Q(
        n1087) );
  AO22X1 U172 ( .IN1(n40), .IN2(n78), .IN3(\mem[30][14] ), .IN4(n1988), .Q(
        n1088) );
  AO22X1 U173 ( .IN1(n41), .IN2(n1928), .IN3(\mem[30][15] ), .IN4(n1988), .Q(
        n1089) );
  AO22X1 U174 ( .IN1(n42), .IN2(n1927), .IN3(\mem[30][16] ), .IN4(n1988), .Q(
        n1090) );
  AO22X1 U175 ( .IN1(n43), .IN2(n78), .IN3(\mem[30][17] ), .IN4(n1988), .Q(
        n1091) );
  AO22X1 U176 ( .IN1(n44), .IN2(n1928), .IN3(\mem[30][18] ), .IN4(n1988), .Q(
        n1092) );
  AO22X1 U177 ( .IN1(n45), .IN2(n1927), .IN3(\mem[30][19] ), .IN4(n1988), .Q(
        n1093) );
  AO22X1 U178 ( .IN1(n46), .IN2(n78), .IN3(\mem[30][20] ), .IN4(n1988), .Q(
        n1094) );
  AO22X1 U179 ( .IN1(n47), .IN2(n1928), .IN3(\mem[30][21] ), .IN4(n1988), .Q(
        n1095) );
  AO22X1 U180 ( .IN1(n48), .IN2(n1927), .IN3(\mem[30][22] ), .IN4(n1988), .Q(
        n1096) );
  AO22X1 U181 ( .IN1(n49), .IN2(n78), .IN3(\mem[30][23] ), .IN4(n1988), .Q(
        n1097) );
  AO22X1 U182 ( .IN1(n1854), .IN2(n1928), .IN3(\mem[30][24] ), .IN4(n1988), 
        .Q(n1098) );
  AO22X1 U183 ( .IN1(n1853), .IN2(n1927), .IN3(\mem[30][25] ), .IN4(n1988), 
        .Q(n1099) );
  AO22X1 U184 ( .IN1(n1852), .IN2(n1928), .IN3(\mem[30][26] ), .IN4(n1987), 
        .Q(n1100) );
  AO22X1 U185 ( .IN1(n1851), .IN2(n1927), .IN3(\mem[30][27] ), .IN4(n1988), 
        .Q(n1101) );
  AO22X1 U186 ( .IN1(n1850), .IN2(n1928), .IN3(\mem[30][28] ), .IN4(n1987), 
        .Q(n1102) );
  AO22X1 U187 ( .IN1(n1849), .IN2(n1927), .IN3(\mem[30][29] ), .IN4(n1988), 
        .Q(n1103) );
  AO22X1 U188 ( .IN1(n1848), .IN2(n1928), .IN3(\mem[30][30] ), .IN4(n1987), 
        .Q(n1104) );
  AO22X1 U189 ( .IN1(n1845), .IN2(n1927), .IN3(\mem[30][31] ), .IN4(n1987), 
        .Q(n1105) );
  AO22X1 U191 ( .IN1(n1844), .IN2(n1926), .IN3(\mem[31][0] ), .IN4(n1985), .Q(
        n1106) );
  AO22X1 U192 ( .IN1(n1843), .IN2(n1925), .IN3(\mem[31][1] ), .IN4(n1985), .Q(
        n1107) );
  AO22X1 U193 ( .IN1(n61), .IN2(n80), .IN3(\mem[31][2] ), .IN4(n1985), .Q(
        n1108) );
  AO22X1 U194 ( .IN1(n62), .IN2(n1926), .IN3(\mem[31][3] ), .IN4(n1985), .Q(
        n1109) );
  AO22X1 U195 ( .IN1(n63), .IN2(n1925), .IN3(\mem[31][4] ), .IN4(n1985), .Q(
        n1110) );
  AO22X1 U196 ( .IN1(n64), .IN2(n80), .IN3(\mem[31][5] ), .IN4(n1985), .Q(
        n1111) );
  AO22X1 U197 ( .IN1(n65), .IN2(n1926), .IN3(\mem[31][6] ), .IN4(n1985), .Q(
        n1112) );
  AO22X1 U198 ( .IN1(n66), .IN2(n1925), .IN3(\mem[31][7] ), .IN4(n1985), .Q(
        n1113) );
  AO22X1 U199 ( .IN1(n67), .IN2(n80), .IN3(\mem[31][8] ), .IN4(n1985), .Q(
        n1114) );
  AO22X1 U200 ( .IN1(n68), .IN2(n1926), .IN3(\mem[31][9] ), .IN4(n1985), .Q(
        n1115) );
  AO22X1 U201 ( .IN1(n69), .IN2(n1925), .IN3(\mem[31][10] ), .IN4(n1985), .Q(
        n1116) );
  AO22X1 U202 ( .IN1(n70), .IN2(n80), .IN3(\mem[31][11] ), .IN4(n1985), .Q(
        n1117) );
  AO22X1 U203 ( .IN1(n71), .IN2(n1926), .IN3(\mem[31][12] ), .IN4(n1986), .Q(
        n1118) );
  AO22X1 U204 ( .IN1(n1876), .IN2(n1925), .IN3(\mem[31][13] ), .IN4(n1986), 
        .Q(n1119) );
  AO22X1 U205 ( .IN1(n1874), .IN2(n80), .IN3(\mem[31][14] ), .IN4(n1986), .Q(
        n1120) );
  AO22X1 U206 ( .IN1(n1872), .IN2(n1926), .IN3(\mem[31][15] ), .IN4(n1986), 
        .Q(n1121) );
  AO22X1 U207 ( .IN1(n1870), .IN2(n1925), .IN3(\mem[31][16] ), .IN4(n1986), 
        .Q(n1122) );
  AO22X1 U208 ( .IN1(n1868), .IN2(n80), .IN3(\mem[31][17] ), .IN4(n1986), .Q(
        n1123) );
  AO22X1 U209 ( .IN1(n1866), .IN2(n1926), .IN3(\mem[31][18] ), .IN4(n1986), 
        .Q(n1124) );
  AO22X1 U210 ( .IN1(n1864), .IN2(n1925), .IN3(\mem[31][19] ), .IN4(n1986), 
        .Q(n1125) );
  AO22X1 U211 ( .IN1(n1862), .IN2(n80), .IN3(\mem[31][20] ), .IN4(n1986), .Q(
        n1126) );
  AO22X1 U212 ( .IN1(n1860), .IN2(n1926), .IN3(\mem[31][21] ), .IN4(n1986), 
        .Q(n1127) );
  AO22X1 U213 ( .IN1(n1858), .IN2(n1925), .IN3(\mem[31][22] ), .IN4(n1986), 
        .Q(n1128) );
  AO22X1 U214 ( .IN1(n1856), .IN2(n80), .IN3(\mem[31][23] ), .IN4(n1986), .Q(
        n1129) );
  AO22X1 U215 ( .IN1(n50), .IN2(n1926), .IN3(\mem[31][24] ), .IN4(n1986), .Q(
        n1130) );
  AO22X1 U216 ( .IN1(n51), .IN2(n1925), .IN3(\mem[31][25] ), .IN4(n1986), .Q(
        n1131) );
  AO22X1 U217 ( .IN1(n52), .IN2(n1926), .IN3(\mem[31][26] ), .IN4(n1985), .Q(
        n1132) );
  AO22X1 U218 ( .IN1(n53), .IN2(n1925), .IN3(\mem[31][27] ), .IN4(n1985), .Q(
        n1133) );
  AO22X1 U219 ( .IN1(n54), .IN2(n1926), .IN3(\mem[31][28] ), .IN4(n1986), .Q(
        n1134) );
  AO22X1 U220 ( .IN1(n55), .IN2(n1925), .IN3(\mem[31][29] ), .IN4(n1985), .Q(
        n1135) );
  AO22X1 U221 ( .IN1(n56), .IN2(n1926), .IN3(\mem[31][30] ), .IN4(n1986), .Q(
        n1136) );
  AO22X1 U222 ( .IN1(n57), .IN2(n1925), .IN3(\mem[31][31] ), .IN4(n1985), .Q(
        n1137) );
  AND2X1 U224 ( .IN1(\mem[0][0] ), .IN2(nrst), .Q(n114) );
  AND2X1 U225 ( .IN1(\mem[0][1] ), .IN2(nrst), .Q(n115) );
  AND2X1 U226 ( .IN1(\mem[0][2] ), .IN2(nrst), .Q(n116) );
  AND2X1 U227 ( .IN1(\mem[0][3] ), .IN2(nrst), .Q(n117) );
  AND2X1 U228 ( .IN1(\mem[0][4] ), .IN2(nrst), .Q(n118) );
  AND2X1 U229 ( .IN1(\mem[0][5] ), .IN2(nrst), .Q(n119) );
  AND2X1 U230 ( .IN1(\mem[0][6] ), .IN2(nrst), .Q(n120) );
  AND2X1 U231 ( .IN1(\mem[0][7] ), .IN2(nrst), .Q(n121) );
  AND2X1 U232 ( .IN1(\mem[0][8] ), .IN2(nrst), .Q(n122) );
  AND2X1 U233 ( .IN1(\mem[0][9] ), .IN2(nrst), .Q(n123) );
  AND2X1 U234 ( .IN1(\mem[0][10] ), .IN2(nrst), .Q(n124) );
  AND2X1 U235 ( .IN1(\mem[0][11] ), .IN2(nrst), .Q(n125) );
  AND2X1 U236 ( .IN1(\mem[0][12] ), .IN2(nrst), .Q(n126) );
  AND2X1 U237 ( .IN1(\mem[0][13] ), .IN2(nrst), .Q(n127) );
  AND2X1 U238 ( .IN1(\mem[0][14] ), .IN2(nrst), .Q(n128) );
  AND2X1 U239 ( .IN1(\mem[0][15] ), .IN2(nrst), .Q(n129) );
  AND2X1 U240 ( .IN1(\mem[0][16] ), .IN2(nrst), .Q(n130) );
  AND2X1 U241 ( .IN1(\mem[0][17] ), .IN2(nrst), .Q(n131) );
  AND2X1 U242 ( .IN1(\mem[0][18] ), .IN2(nrst), .Q(n132) );
  AND2X1 U243 ( .IN1(\mem[0][19] ), .IN2(nrst), .Q(n133) );
  AND2X1 U244 ( .IN1(\mem[0][20] ), .IN2(nrst), .Q(n134) );
  AND2X1 U245 ( .IN1(\mem[0][21] ), .IN2(nrst), .Q(n135) );
  AND2X1 U246 ( .IN1(\mem[0][22] ), .IN2(nrst), .Q(n136) );
  AND2X1 U247 ( .IN1(\mem[0][23] ), .IN2(nrst), .Q(n137) );
  AND2X1 U248 ( .IN1(\mem[0][24] ), .IN2(nrst), .Q(n138) );
  AND2X1 U249 ( .IN1(\mem[0][25] ), .IN2(nrst), .Q(n139) );
  AND2X1 U250 ( .IN1(\mem[0][26] ), .IN2(nrst), .Q(n140) );
  AND2X1 U251 ( .IN1(\mem[0][27] ), .IN2(nrst), .Q(n141) );
  AND2X1 U252 ( .IN1(\mem[0][28] ), .IN2(nrst), .Q(n142) );
  AND2X1 U253 ( .IN1(\mem[0][29] ), .IN2(nrst), .Q(n143) );
  AND2X1 U254 ( .IN1(\mem[0][30] ), .IN2(nrst), .Q(n144) );
  AND2X1 U255 ( .IN1(\mem[0][31] ), .IN2(nrst), .Q(n145) );
  AO22X1 U256 ( .IN1(n58), .IN2(n1924), .IN3(\mem[1][0] ), .IN4(n1983), .Q(
        n146) );
  AO22X1 U257 ( .IN1(n60), .IN2(n1923), .IN3(\mem[1][1] ), .IN4(n1983), .Q(
        n147) );
  AO22X1 U258 ( .IN1(n61), .IN2(n82), .IN3(\mem[1][2] ), .IN4(n1983), .Q(n148)
         );
  AO22X1 U259 ( .IN1(n62), .IN2(n1924), .IN3(\mem[1][3] ), .IN4(n1983), .Q(
        n149) );
  AO22X1 U260 ( .IN1(n63), .IN2(n1923), .IN3(\mem[1][4] ), .IN4(n1983), .Q(
        n150) );
  AO22X1 U261 ( .IN1(n64), .IN2(n82), .IN3(\mem[1][5] ), .IN4(n1983), .Q(n151)
         );
  AO22X1 U262 ( .IN1(n65), .IN2(n1924), .IN3(\mem[1][6] ), .IN4(n1983), .Q(
        n152) );
  AO22X1 U263 ( .IN1(n66), .IN2(n1923), .IN3(\mem[1][7] ), .IN4(n1983), .Q(
        n153) );
  AO22X1 U264 ( .IN1(n67), .IN2(n82), .IN3(\mem[1][8] ), .IN4(n1983), .Q(n154)
         );
  AO22X1 U265 ( .IN1(n68), .IN2(n1924), .IN3(\mem[1][9] ), .IN4(n1983), .Q(
        n155) );
  AO22X1 U266 ( .IN1(n69), .IN2(n1923), .IN3(\mem[1][10] ), .IN4(n1983), .Q(
        n156) );
  AO22X1 U267 ( .IN1(n70), .IN2(n82), .IN3(\mem[1][11] ), .IN4(n1983), .Q(n157) );
  AO22X1 U268 ( .IN1(n71), .IN2(n1924), .IN3(\mem[1][12] ), .IN4(n1984), .Q(
        n158) );
  AO22X1 U269 ( .IN1(n1875), .IN2(n1923), .IN3(\mem[1][13] ), .IN4(n1984), .Q(
        n159) );
  AO22X1 U270 ( .IN1(n1873), .IN2(n82), .IN3(\mem[1][14] ), .IN4(n1984), .Q(
        n160) );
  AO22X1 U271 ( .IN1(n1871), .IN2(n1924), .IN3(\mem[1][15] ), .IN4(n1984), .Q(
        n161) );
  AO22X1 U272 ( .IN1(n1869), .IN2(n1923), .IN3(\mem[1][16] ), .IN4(n1984), .Q(
        n162) );
  AO22X1 U273 ( .IN1(n1867), .IN2(n82), .IN3(\mem[1][17] ), .IN4(n1984), .Q(
        n163) );
  AO22X1 U274 ( .IN1(n1865), .IN2(n1924), .IN3(\mem[1][18] ), .IN4(n1984), .Q(
        n164) );
  AO22X1 U275 ( .IN1(n1863), .IN2(n1923), .IN3(\mem[1][19] ), .IN4(n1984), .Q(
        n165) );
  AO22X1 U276 ( .IN1(n1861), .IN2(n82), .IN3(\mem[1][20] ), .IN4(n1984), .Q(
        n166) );
  AO22X1 U277 ( .IN1(n1859), .IN2(n1924), .IN3(\mem[1][21] ), .IN4(n1984), .Q(
        n167) );
  AO22X1 U278 ( .IN1(n1857), .IN2(n1923), .IN3(\mem[1][22] ), .IN4(n1984), .Q(
        n168) );
  AO22X1 U279 ( .IN1(n1855), .IN2(n82), .IN3(\mem[1][23] ), .IN4(n1984), .Q(
        n169) );
  AO22X1 U280 ( .IN1(n1854), .IN2(n1924), .IN3(\mem[1][24] ), .IN4(n1984), .Q(
        n170) );
  AO22X1 U281 ( .IN1(n1853), .IN2(n1923), .IN3(\mem[1][25] ), .IN4(n1984), .Q(
        n171) );
  AO22X1 U282 ( .IN1(n1852), .IN2(n1924), .IN3(\mem[1][26] ), .IN4(n1983), .Q(
        n172) );
  AO22X1 U283 ( .IN1(n1851), .IN2(n1923), .IN3(\mem[1][27] ), .IN4(n1984), .Q(
        n173) );
  AO22X1 U284 ( .IN1(n1850), .IN2(n1924), .IN3(\mem[1][28] ), .IN4(n1983), .Q(
        n174) );
  AO22X1 U285 ( .IN1(n1849), .IN2(n1923), .IN3(\mem[1][29] ), .IN4(n1984), .Q(
        n175) );
  AO22X1 U286 ( .IN1(n1848), .IN2(n1924), .IN3(\mem[1][30] ), .IN4(n1983), .Q(
        n176) );
  AO22X1 U287 ( .IN1(n1845), .IN2(n1923), .IN3(\mem[1][31] ), .IN4(n1983), .Q(
        n177) );
  AO22X1 U289 ( .IN1(n1844), .IN2(n1922), .IN3(\mem[2][0] ), .IN4(n1981), .Q(
        n178) );
  AO22X1 U290 ( .IN1(n1843), .IN2(n1921), .IN3(\mem[2][1] ), .IN4(n1981), .Q(
        n179) );
  AO22X1 U291 ( .IN1(n61), .IN2(n85), .IN3(\mem[2][2] ), .IN4(n1981), .Q(n180)
         );
  AO22X1 U292 ( .IN1(n62), .IN2(n1922), .IN3(\mem[2][3] ), .IN4(n1981), .Q(
        n181) );
  AO22X1 U293 ( .IN1(n63), .IN2(n1921), .IN3(\mem[2][4] ), .IN4(n1981), .Q(
        n182) );
  AO22X1 U294 ( .IN1(n64), .IN2(n85), .IN3(\mem[2][5] ), .IN4(n1981), .Q(n183)
         );
  AO22X1 U295 ( .IN1(n65), .IN2(n1922), .IN3(\mem[2][6] ), .IN4(n1981), .Q(
        n184) );
  AO22X1 U296 ( .IN1(n66), .IN2(n1921), .IN3(\mem[2][7] ), .IN4(n1981), .Q(
        n185) );
  AO22X1 U297 ( .IN1(n67), .IN2(n85), .IN3(\mem[2][8] ), .IN4(n1981), .Q(n186)
         );
  AO22X1 U298 ( .IN1(n68), .IN2(n1922), .IN3(\mem[2][9] ), .IN4(n1981), .Q(
        n187) );
  AO22X1 U299 ( .IN1(n69), .IN2(n1921), .IN3(\mem[2][10] ), .IN4(n1981), .Q(
        n188) );
  AO22X1 U300 ( .IN1(n70), .IN2(n85), .IN3(\mem[2][11] ), .IN4(n1981), .Q(n189) );
  AO22X1 U301 ( .IN1(n71), .IN2(n1922), .IN3(\mem[2][12] ), .IN4(n1982), .Q(
        n190) );
  AO22X1 U302 ( .IN1(n38), .IN2(n1921), .IN3(\mem[2][13] ), .IN4(n1982), .Q(
        n191) );
  AO22X1 U303 ( .IN1(n40), .IN2(n85), .IN3(\mem[2][14] ), .IN4(n1982), .Q(n192) );
  AO22X1 U304 ( .IN1(n41), .IN2(n1922), .IN3(\mem[2][15] ), .IN4(n1982), .Q(
        n193) );
  AO22X1 U305 ( .IN1(n42), .IN2(n1921), .IN3(\mem[2][16] ), .IN4(n1982), .Q(
        n194) );
  AO22X1 U306 ( .IN1(n43), .IN2(n85), .IN3(\mem[2][17] ), .IN4(n1982), .Q(n195) );
  AO22X1 U307 ( .IN1(n44), .IN2(n1922), .IN3(\mem[2][18] ), .IN4(n1982), .Q(
        n196) );
  AO22X1 U308 ( .IN1(n45), .IN2(n1921), .IN3(\mem[2][19] ), .IN4(n1982), .Q(
        n197) );
  AO22X1 U309 ( .IN1(n46), .IN2(n85), .IN3(\mem[2][20] ), .IN4(n1982), .Q(n198) );
  AO22X1 U310 ( .IN1(n47), .IN2(n1922), .IN3(\mem[2][21] ), .IN4(n1982), .Q(
        n199) );
  AO22X1 U311 ( .IN1(n48), .IN2(n1921), .IN3(\mem[2][22] ), .IN4(n1982), .Q(
        n200) );
  AO22X1 U312 ( .IN1(n49), .IN2(n85), .IN3(\mem[2][23] ), .IN4(n1982), .Q(n201) );
  AO22X1 U313 ( .IN1(n50), .IN2(n1922), .IN3(\mem[2][24] ), .IN4(n1982), .Q(
        n202) );
  AO22X1 U314 ( .IN1(n51), .IN2(n1921), .IN3(\mem[2][25] ), .IN4(n1982), .Q(
        n203) );
  AO22X1 U315 ( .IN1(n52), .IN2(n1922), .IN3(\mem[2][26] ), .IN4(n1981), .Q(
        n204) );
  AO22X1 U316 ( .IN1(n53), .IN2(n1921), .IN3(\mem[2][27] ), .IN4(n1981), .Q(
        n205) );
  AO22X1 U317 ( .IN1(n54), .IN2(n1922), .IN3(\mem[2][28] ), .IN4(n1982), .Q(
        n206) );
  AO22X1 U318 ( .IN1(n55), .IN2(n1921), .IN3(\mem[2][29] ), .IN4(n1981), .Q(
        n207) );
  AO22X1 U319 ( .IN1(n56), .IN2(n1922), .IN3(\mem[2][30] ), .IN4(n1982), .Q(
        n208) );
  AO22X1 U320 ( .IN1(n57), .IN2(n1921), .IN3(\mem[2][31] ), .IN4(n1981), .Q(
        n209) );
  AO22X1 U322 ( .IN1(n58), .IN2(n1920), .IN3(\mem[3][0] ), .IN4(n1979), .Q(
        n210) );
  AO22X1 U323 ( .IN1(n60), .IN2(n1919), .IN3(\mem[3][1] ), .IN4(n1979), .Q(
        n211) );
  AO22X1 U324 ( .IN1(n61), .IN2(n87), .IN3(\mem[3][2] ), .IN4(n1979), .Q(n212)
         );
  AO22X1 U325 ( .IN1(n62), .IN2(n1920), .IN3(\mem[3][3] ), .IN4(n1979), .Q(
        n213) );
  AO22X1 U326 ( .IN1(n63), .IN2(n1919), .IN3(\mem[3][4] ), .IN4(n1979), .Q(
        n214) );
  AO22X1 U327 ( .IN1(n64), .IN2(n87), .IN3(\mem[3][5] ), .IN4(n1979), .Q(n215)
         );
  AO22X1 U328 ( .IN1(n65), .IN2(n1920), .IN3(\mem[3][6] ), .IN4(n1979), .Q(
        n216) );
  AO22X1 U329 ( .IN1(n66), .IN2(n1919), .IN3(\mem[3][7] ), .IN4(n1979), .Q(
        n217) );
  AO22X1 U330 ( .IN1(n67), .IN2(n87), .IN3(\mem[3][8] ), .IN4(n1979), .Q(n218)
         );
  AO22X1 U331 ( .IN1(n68), .IN2(n1920), .IN3(\mem[3][9] ), .IN4(n1979), .Q(
        n219) );
  AO22X1 U332 ( .IN1(n69), .IN2(n1919), .IN3(\mem[3][10] ), .IN4(n1979), .Q(
        n220) );
  AO22X1 U333 ( .IN1(n70), .IN2(n87), .IN3(\mem[3][11] ), .IN4(n1979), .Q(n221) );
  AO22X1 U334 ( .IN1(n71), .IN2(n1920), .IN3(\mem[3][12] ), .IN4(n1980), .Q(
        n222) );
  AO22X1 U335 ( .IN1(n1876), .IN2(n1919), .IN3(\mem[3][13] ), .IN4(n1980), .Q(
        n223) );
  AO22X1 U336 ( .IN1(n1874), .IN2(n87), .IN3(\mem[3][14] ), .IN4(n1980), .Q(
        n224) );
  AO22X1 U337 ( .IN1(n1872), .IN2(n1920), .IN3(\mem[3][15] ), .IN4(n1980), .Q(
        n225) );
  AO22X1 U338 ( .IN1(n1870), .IN2(n1919), .IN3(\mem[3][16] ), .IN4(n1980), .Q(
        n226) );
  AO22X1 U339 ( .IN1(n1868), .IN2(n87), .IN3(\mem[3][17] ), .IN4(n1980), .Q(
        n227) );
  AO22X1 U340 ( .IN1(n1866), .IN2(n1920), .IN3(\mem[3][18] ), .IN4(n1980), .Q(
        n228) );
  AO22X1 U341 ( .IN1(n1864), .IN2(n1919), .IN3(\mem[3][19] ), .IN4(n1980), .Q(
        n229) );
  AO22X1 U342 ( .IN1(n1862), .IN2(n87), .IN3(\mem[3][20] ), .IN4(n1980), .Q(
        n230) );
  AO22X1 U343 ( .IN1(n1860), .IN2(n1920), .IN3(\mem[3][21] ), .IN4(n1980), .Q(
        n231) );
  AO22X1 U344 ( .IN1(n1858), .IN2(n1919), .IN3(\mem[3][22] ), .IN4(n1980), .Q(
        n232) );
  AO22X1 U345 ( .IN1(n1856), .IN2(n87), .IN3(\mem[3][23] ), .IN4(n1980), .Q(
        n233) );
  AO22X1 U346 ( .IN1(n1854), .IN2(n1920), .IN3(\mem[3][24] ), .IN4(n1980), .Q(
        n234) );
  AO22X1 U347 ( .IN1(n1853), .IN2(n1919), .IN3(\mem[3][25] ), .IN4(n1980), .Q(
        n235) );
  AO22X1 U348 ( .IN1(n1852), .IN2(n1920), .IN3(\mem[3][26] ), .IN4(n1979), .Q(
        n236) );
  AO22X1 U349 ( .IN1(n1851), .IN2(n1919), .IN3(\mem[3][27] ), .IN4(n1980), .Q(
        n237) );
  AO22X1 U350 ( .IN1(n1850), .IN2(n1920), .IN3(\mem[3][28] ), .IN4(n1979), .Q(
        n238) );
  AO22X1 U351 ( .IN1(n1849), .IN2(n1919), .IN3(\mem[3][29] ), .IN4(n1980), .Q(
        n239) );
  AO22X1 U352 ( .IN1(n1848), .IN2(n1920), .IN3(\mem[3][30] ), .IN4(n1979), .Q(
        n240) );
  AO22X1 U353 ( .IN1(n1845), .IN2(n1919), .IN3(\mem[3][31] ), .IN4(n1979), .Q(
        n241) );
  AO22X1 U355 ( .IN1(n1844), .IN2(n1918), .IN3(\mem[4][0] ), .IN4(n1977), .Q(
        n242) );
  AO22X1 U356 ( .IN1(n1843), .IN2(n1917), .IN3(\mem[4][1] ), .IN4(n1977), .Q(
        n243) );
  AO22X1 U357 ( .IN1(n61), .IN2(n88), .IN3(\mem[4][2] ), .IN4(n1977), .Q(n244)
         );
  AO22X1 U358 ( .IN1(n62), .IN2(n1918), .IN3(\mem[4][3] ), .IN4(n1977), .Q(
        n245) );
  AO22X1 U359 ( .IN1(n63), .IN2(n1917), .IN3(\mem[4][4] ), .IN4(n1977), .Q(
        n246) );
  AO22X1 U360 ( .IN1(n64), .IN2(n88), .IN3(\mem[4][5] ), .IN4(n1977), .Q(n247)
         );
  AO22X1 U361 ( .IN1(n65), .IN2(n1918), .IN3(\mem[4][6] ), .IN4(n1977), .Q(
        n248) );
  AO22X1 U362 ( .IN1(n66), .IN2(n1917), .IN3(\mem[4][7] ), .IN4(n1977), .Q(
        n249) );
  AO22X1 U363 ( .IN1(n67), .IN2(n88), .IN3(\mem[4][8] ), .IN4(n1977), .Q(n250)
         );
  AO22X1 U364 ( .IN1(n68), .IN2(n1918), .IN3(\mem[4][9] ), .IN4(n1977), .Q(
        n251) );
  AO22X1 U365 ( .IN1(n69), .IN2(n1917), .IN3(\mem[4][10] ), .IN4(n1977), .Q(
        n252) );
  AO22X1 U366 ( .IN1(n70), .IN2(n88), .IN3(\mem[4][11] ), .IN4(n1977), .Q(n253) );
  AO22X1 U367 ( .IN1(n71), .IN2(n1918), .IN3(\mem[4][12] ), .IN4(n1978), .Q(
        n254) );
  AO22X1 U368 ( .IN1(n1875), .IN2(n1917), .IN3(\mem[4][13] ), .IN4(n1978), .Q(
        n255) );
  AO22X1 U369 ( .IN1(n1873), .IN2(n88), .IN3(\mem[4][14] ), .IN4(n1978), .Q(
        n256) );
  AO22X1 U370 ( .IN1(n1871), .IN2(n1918), .IN3(\mem[4][15] ), .IN4(n1978), .Q(
        n257) );
  AO22X1 U371 ( .IN1(n1869), .IN2(n1917), .IN3(\mem[4][16] ), .IN4(n1978), .Q(
        n258) );
  AO22X1 U372 ( .IN1(n1867), .IN2(n88), .IN3(\mem[4][17] ), .IN4(n1978), .Q(
        n259) );
  AO22X1 U373 ( .IN1(n1865), .IN2(n1918), .IN3(\mem[4][18] ), .IN4(n1978), .Q(
        n260) );
  AO22X1 U374 ( .IN1(n1863), .IN2(n1917), .IN3(\mem[4][19] ), .IN4(n1978), .Q(
        n261) );
  AO22X1 U375 ( .IN1(n1861), .IN2(n88), .IN3(\mem[4][20] ), .IN4(n1978), .Q(
        n262) );
  AO22X1 U376 ( .IN1(n1859), .IN2(n1918), .IN3(\mem[4][21] ), .IN4(n1978), .Q(
        n263) );
  AO22X1 U377 ( .IN1(n1857), .IN2(n1917), .IN3(\mem[4][22] ), .IN4(n1978), .Q(
        n264) );
  AO22X1 U378 ( .IN1(n1855), .IN2(n88), .IN3(\mem[4][23] ), .IN4(n1978), .Q(
        n265) );
  AO22X1 U379 ( .IN1(n50), .IN2(n1918), .IN3(\mem[4][24] ), .IN4(n1978), .Q(
        n266) );
  AO22X1 U380 ( .IN1(n51), .IN2(n1917), .IN3(\mem[4][25] ), .IN4(n1978), .Q(
        n267) );
  AO22X1 U381 ( .IN1(n52), .IN2(n1918), .IN3(\mem[4][26] ), .IN4(n1977), .Q(
        n268) );
  AO22X1 U382 ( .IN1(n53), .IN2(n1917), .IN3(\mem[4][27] ), .IN4(n1977), .Q(
        n269) );
  AO22X1 U383 ( .IN1(n54), .IN2(n1918), .IN3(\mem[4][28] ), .IN4(n1978), .Q(
        n270) );
  AO22X1 U384 ( .IN1(n55), .IN2(n1917), .IN3(\mem[4][29] ), .IN4(n1977), .Q(
        n271) );
  AO22X1 U385 ( .IN1(n56), .IN2(n1918), .IN3(\mem[4][30] ), .IN4(n1978), .Q(
        n272) );
  AO22X1 U386 ( .IN1(n57), .IN2(n1917), .IN3(\mem[4][31] ), .IN4(n1977), .Q(
        n273) );
  AO22X1 U388 ( .IN1(n58), .IN2(n1916), .IN3(\mem[5][0] ), .IN4(n1975), .Q(
        n274) );
  AO22X1 U389 ( .IN1(n60), .IN2(n1915), .IN3(\mem[5][1] ), .IN4(n1975), .Q(
        n275) );
  AO22X1 U390 ( .IN1(n61), .IN2(n89), .IN3(\mem[5][2] ), .IN4(n1975), .Q(n276)
         );
  AO22X1 U391 ( .IN1(n62), .IN2(n1916), .IN3(\mem[5][3] ), .IN4(n1975), .Q(
        n277) );
  AO22X1 U392 ( .IN1(n63), .IN2(n1915), .IN3(\mem[5][4] ), .IN4(n1975), .Q(
        n278) );
  AO22X1 U393 ( .IN1(n64), .IN2(n89), .IN3(\mem[5][5] ), .IN4(n1975), .Q(n279)
         );
  AO22X1 U394 ( .IN1(n65), .IN2(n1916), .IN3(\mem[5][6] ), .IN4(n1975), .Q(
        n280) );
  AO22X1 U395 ( .IN1(n66), .IN2(n1915), .IN3(\mem[5][7] ), .IN4(n1975), .Q(
        n281) );
  AO22X1 U396 ( .IN1(n67), .IN2(n89), .IN3(\mem[5][8] ), .IN4(n1975), .Q(n282)
         );
  AO22X1 U397 ( .IN1(n68), .IN2(n1916), .IN3(\mem[5][9] ), .IN4(n1975), .Q(
        n283) );
  AO22X1 U398 ( .IN1(n69), .IN2(n1915), .IN3(\mem[5][10] ), .IN4(n1975), .Q(
        n284) );
  AO22X1 U399 ( .IN1(n70), .IN2(n89), .IN3(\mem[5][11] ), .IN4(n1975), .Q(n285) );
  AO22X1 U400 ( .IN1(n71), .IN2(n1916), .IN3(\mem[5][12] ), .IN4(n1976), .Q(
        n286) );
  AO22X1 U401 ( .IN1(n38), .IN2(n1915), .IN3(\mem[5][13] ), .IN4(n1976), .Q(
        n287) );
  AO22X1 U402 ( .IN1(n40), .IN2(n89), .IN3(\mem[5][14] ), .IN4(n1976), .Q(n288) );
  AO22X1 U403 ( .IN1(n41), .IN2(n1916), .IN3(\mem[5][15] ), .IN4(n1976), .Q(
        n289) );
  AO22X1 U404 ( .IN1(n42), .IN2(n1915), .IN3(\mem[5][16] ), .IN4(n1976), .Q(
        n290) );
  AO22X1 U405 ( .IN1(n43), .IN2(n89), .IN3(\mem[5][17] ), .IN4(n1976), .Q(n291) );
  AO22X1 U406 ( .IN1(n44), .IN2(n1916), .IN3(\mem[5][18] ), .IN4(n1976), .Q(
        n292) );
  AO22X1 U407 ( .IN1(n45), .IN2(n1915), .IN3(\mem[5][19] ), .IN4(n1976), .Q(
        n293) );
  AO22X1 U408 ( .IN1(n46), .IN2(n89), .IN3(\mem[5][20] ), .IN4(n1976), .Q(n294) );
  AO22X1 U409 ( .IN1(n47), .IN2(n1916), .IN3(\mem[5][21] ), .IN4(n1976), .Q(
        n295) );
  AO22X1 U410 ( .IN1(n48), .IN2(n1915), .IN3(\mem[5][22] ), .IN4(n1976), .Q(
        n296) );
  AO22X1 U411 ( .IN1(n49), .IN2(n89), .IN3(\mem[5][23] ), .IN4(n1976), .Q(n297) );
  AO22X1 U412 ( .IN1(n1854), .IN2(n1916), .IN3(\mem[5][24] ), .IN4(n1976), .Q(
        n298) );
  AO22X1 U413 ( .IN1(n1853), .IN2(n1915), .IN3(\mem[5][25] ), .IN4(n1976), .Q(
        n299) );
  AO22X1 U414 ( .IN1(n1852), .IN2(n1916), .IN3(\mem[5][26] ), .IN4(n1975), .Q(
        n300) );
  AO22X1 U415 ( .IN1(n1851), .IN2(n1915), .IN3(\mem[5][27] ), .IN4(n1976), .Q(
        n301) );
  AO22X1 U416 ( .IN1(n1850), .IN2(n1916), .IN3(\mem[5][28] ), .IN4(n1975), .Q(
        n302) );
  AO22X1 U417 ( .IN1(n1849), .IN2(n1915), .IN3(\mem[5][29] ), .IN4(n1976), .Q(
        n303) );
  AO22X1 U418 ( .IN1(n1848), .IN2(n1916), .IN3(\mem[5][30] ), .IN4(n1975), .Q(
        n304) );
  AO22X1 U419 ( .IN1(n1845), .IN2(n1915), .IN3(\mem[5][31] ), .IN4(n1975), .Q(
        n305) );
  AO22X1 U421 ( .IN1(n1844), .IN2(n1914), .IN3(\mem[6][0] ), .IN4(n1973), .Q(
        n306) );
  AO22X1 U422 ( .IN1(n1843), .IN2(n1913), .IN3(\mem[6][1] ), .IN4(n1973), .Q(
        n307) );
  AO22X1 U423 ( .IN1(n61), .IN2(n90), .IN3(\mem[6][2] ), .IN4(n1973), .Q(n308)
         );
  AO22X1 U424 ( .IN1(n62), .IN2(n1914), .IN3(\mem[6][3] ), .IN4(n1973), .Q(
        n309) );
  AO22X1 U425 ( .IN1(n63), .IN2(n1913), .IN3(\mem[6][4] ), .IN4(n1973), .Q(
        n310) );
  AO22X1 U426 ( .IN1(n64), .IN2(n90), .IN3(\mem[6][5] ), .IN4(n1973), .Q(n311)
         );
  AO22X1 U427 ( .IN1(n65), .IN2(n1914), .IN3(\mem[6][6] ), .IN4(n1973), .Q(
        n312) );
  AO22X1 U428 ( .IN1(n66), .IN2(n1913), .IN3(\mem[6][7] ), .IN4(n1973), .Q(
        n313) );
  AO22X1 U429 ( .IN1(n67), .IN2(n90), .IN3(\mem[6][8] ), .IN4(n1973), .Q(n314)
         );
  AO22X1 U430 ( .IN1(n68), .IN2(n1914), .IN3(\mem[6][9] ), .IN4(n1973), .Q(
        n315) );
  AO22X1 U431 ( .IN1(n69), .IN2(n1913), .IN3(\mem[6][10] ), .IN4(n1973), .Q(
        n316) );
  AO22X1 U432 ( .IN1(n70), .IN2(n90), .IN3(\mem[6][11] ), .IN4(n1973), .Q(n317) );
  AO22X1 U433 ( .IN1(n71), .IN2(n1914), .IN3(\mem[6][12] ), .IN4(n1974), .Q(
        n318) );
  AO22X1 U434 ( .IN1(n1876), .IN2(n1913), .IN3(\mem[6][13] ), .IN4(n1974), .Q(
        n319) );
  AO22X1 U435 ( .IN1(n1874), .IN2(n90), .IN3(\mem[6][14] ), .IN4(n1974), .Q(
        n320) );
  AO22X1 U436 ( .IN1(n1872), .IN2(n1914), .IN3(\mem[6][15] ), .IN4(n1974), .Q(
        n321) );
  AO22X1 U437 ( .IN1(n1870), .IN2(n1913), .IN3(\mem[6][16] ), .IN4(n1974), .Q(
        n322) );
  AO22X1 U438 ( .IN1(n1868), .IN2(n90), .IN3(\mem[6][17] ), .IN4(n1974), .Q(
        n323) );
  AO22X1 U439 ( .IN1(n1866), .IN2(n1914), .IN3(\mem[6][18] ), .IN4(n1974), .Q(
        n324) );
  AO22X1 U440 ( .IN1(n1864), .IN2(n1913), .IN3(\mem[6][19] ), .IN4(n1974), .Q(
        n325) );
  AO22X1 U441 ( .IN1(n1862), .IN2(n90), .IN3(\mem[6][20] ), .IN4(n1974), .Q(
        n326) );
  AO22X1 U442 ( .IN1(n1860), .IN2(n1914), .IN3(\mem[6][21] ), .IN4(n1974), .Q(
        n327) );
  AO22X1 U443 ( .IN1(n1858), .IN2(n1913), .IN3(\mem[6][22] ), .IN4(n1974), .Q(
        n328) );
  AO22X1 U444 ( .IN1(n1856), .IN2(n90), .IN3(\mem[6][23] ), .IN4(n1974), .Q(
        n329) );
  AO22X1 U445 ( .IN1(n50), .IN2(n1914), .IN3(\mem[6][24] ), .IN4(n1974), .Q(
        n330) );
  AO22X1 U446 ( .IN1(n51), .IN2(n1913), .IN3(\mem[6][25] ), .IN4(n1974), .Q(
        n331) );
  AO22X1 U447 ( .IN1(n52), .IN2(n1914), .IN3(\mem[6][26] ), .IN4(n1973), .Q(
        n332) );
  AO22X1 U448 ( .IN1(n53), .IN2(n1913), .IN3(\mem[6][27] ), .IN4(n1973), .Q(
        n333) );
  AO22X1 U449 ( .IN1(n54), .IN2(n1914), .IN3(\mem[6][28] ), .IN4(n1974), .Q(
        n334) );
  AO22X1 U450 ( .IN1(n55), .IN2(n1913), .IN3(\mem[6][29] ), .IN4(n1973), .Q(
        n335) );
  AO22X1 U451 ( .IN1(n56), .IN2(n1914), .IN3(\mem[6][30] ), .IN4(n1974), .Q(
        n336) );
  AO22X1 U452 ( .IN1(n57), .IN2(n1913), .IN3(\mem[6][31] ), .IN4(n1973), .Q(
        n337) );
  AO21X1 U453 ( .IN1(n84), .IN2(n79), .IN3(n1997), .Q(n90) );
  AO22X1 U454 ( .IN1(n58), .IN2(n1912), .IN3(\mem[7][0] ), .IN4(n1971), .Q(
        n338) );
  AO22X1 U455 ( .IN1(n60), .IN2(n1911), .IN3(\mem[7][1] ), .IN4(n1971), .Q(
        n339) );
  AO22X1 U456 ( .IN1(n61), .IN2(n91), .IN3(\mem[7][2] ), .IN4(n1971), .Q(n340)
         );
  AO22X1 U457 ( .IN1(n62), .IN2(n1912), .IN3(\mem[7][3] ), .IN4(n1971), .Q(
        n341) );
  AO22X1 U458 ( .IN1(n63), .IN2(n1911), .IN3(\mem[7][4] ), .IN4(n1971), .Q(
        n342) );
  AO22X1 U459 ( .IN1(n64), .IN2(n91), .IN3(\mem[7][5] ), .IN4(n1971), .Q(n343)
         );
  AO22X1 U460 ( .IN1(n65), .IN2(n1912), .IN3(\mem[7][6] ), .IN4(n1971), .Q(
        n344) );
  AO22X1 U461 ( .IN1(n66), .IN2(n1911), .IN3(\mem[7][7] ), .IN4(n1971), .Q(
        n345) );
  AO22X1 U462 ( .IN1(n67), .IN2(n91), .IN3(\mem[7][8] ), .IN4(n1971), .Q(n346)
         );
  AO22X1 U463 ( .IN1(n68), .IN2(n1912), .IN3(\mem[7][9] ), .IN4(n1971), .Q(
        n347) );
  AO22X1 U464 ( .IN1(n69), .IN2(n1911), .IN3(\mem[7][10] ), .IN4(n1971), .Q(
        n348) );
  AO22X1 U465 ( .IN1(n70), .IN2(n91), .IN3(\mem[7][11] ), .IN4(n1971), .Q(n349) );
  AO22X1 U466 ( .IN1(n71), .IN2(n1912), .IN3(\mem[7][12] ), .IN4(n1972), .Q(
        n350) );
  AO22X1 U467 ( .IN1(n1875), .IN2(n1911), .IN3(\mem[7][13] ), .IN4(n1972), .Q(
        n351) );
  AO22X1 U468 ( .IN1(n1873), .IN2(n91), .IN3(\mem[7][14] ), .IN4(n1972), .Q(
        n352) );
  AO22X1 U469 ( .IN1(n1871), .IN2(n1912), .IN3(\mem[7][15] ), .IN4(n1972), .Q(
        n353) );
  AO22X1 U470 ( .IN1(n1869), .IN2(n1911), .IN3(\mem[7][16] ), .IN4(n1972), .Q(
        n354) );
  AO22X1 U471 ( .IN1(n1867), .IN2(n91), .IN3(\mem[7][17] ), .IN4(n1972), .Q(
        n355) );
  AO22X1 U472 ( .IN1(n1865), .IN2(n1912), .IN3(\mem[7][18] ), .IN4(n1972), .Q(
        n356) );
  AO22X1 U473 ( .IN1(n1863), .IN2(n1911), .IN3(\mem[7][19] ), .IN4(n1972), .Q(
        n357) );
  AO22X1 U474 ( .IN1(n1861), .IN2(n91), .IN3(\mem[7][20] ), .IN4(n1972), .Q(
        n358) );
  AO22X1 U475 ( .IN1(n1859), .IN2(n1912), .IN3(\mem[7][21] ), .IN4(n1972), .Q(
        n359) );
  AO22X1 U476 ( .IN1(n1857), .IN2(n1911), .IN3(\mem[7][22] ), .IN4(n1972), .Q(
        n360) );
  AO22X1 U477 ( .IN1(n1855), .IN2(n91), .IN3(\mem[7][23] ), .IN4(n1972), .Q(
        n361) );
  AO22X1 U478 ( .IN1(n1854), .IN2(n1912), .IN3(\mem[7][24] ), .IN4(n1972), .Q(
        n362) );
  AO22X1 U479 ( .IN1(n1853), .IN2(n1911), .IN3(\mem[7][25] ), .IN4(n1972), .Q(
        n363) );
  AO22X1 U480 ( .IN1(n1852), .IN2(n1912), .IN3(\mem[7][26] ), .IN4(n1971), .Q(
        n364) );
  AO22X1 U481 ( .IN1(n1851), .IN2(n1911), .IN3(\mem[7][27] ), .IN4(n1972), .Q(
        n365) );
  AO22X1 U482 ( .IN1(n1850), .IN2(n1912), .IN3(\mem[7][28] ), .IN4(n1971), .Q(
        n366) );
  AO22X1 U483 ( .IN1(n1849), .IN2(n1911), .IN3(\mem[7][29] ), .IN4(n1972), .Q(
        n367) );
  AO22X1 U484 ( .IN1(n1848), .IN2(n1912), .IN3(\mem[7][30] ), .IN4(n1971), .Q(
        n368) );
  AO22X1 U485 ( .IN1(n1845), .IN2(n1911), .IN3(\mem[7][31] ), .IN4(n1971), .Q(
        n369) );
  AO21X1 U486 ( .IN1(n84), .IN2(n81), .IN3(n1997), .Q(n91) );
  AND3X1 U487 ( .IN1(n2001), .IN2(n2000), .IN3(n1837), .Q(n84) );
  AO22X1 U488 ( .IN1(n1844), .IN2(n1910), .IN3(\mem[8][0] ), .IN4(n1969), .Q(
        n370) );
  AO22X1 U489 ( .IN1(n1843), .IN2(n1909), .IN3(\mem[8][1] ), .IN4(n1969), .Q(
        n371) );
  AO22X1 U490 ( .IN1(n61), .IN2(n93), .IN3(\mem[8][2] ), .IN4(n1969), .Q(n372)
         );
  AO22X1 U491 ( .IN1(n62), .IN2(n1910), .IN3(\mem[8][3] ), .IN4(n1969), .Q(
        n373) );
  AO22X1 U492 ( .IN1(n63), .IN2(n1909), .IN3(\mem[8][4] ), .IN4(n1969), .Q(
        n374) );
  AO22X1 U493 ( .IN1(n64), .IN2(n93), .IN3(\mem[8][5] ), .IN4(n1969), .Q(n375)
         );
  AO22X1 U494 ( .IN1(n65), .IN2(n1910), .IN3(\mem[8][6] ), .IN4(n1969), .Q(
        n376) );
  AO22X1 U495 ( .IN1(n66), .IN2(n1909), .IN3(\mem[8][7] ), .IN4(n1969), .Q(
        n377) );
  AO22X1 U496 ( .IN1(n67), .IN2(n93), .IN3(\mem[8][8] ), .IN4(n1969), .Q(n378)
         );
  AO22X1 U497 ( .IN1(n68), .IN2(n1910), .IN3(\mem[8][9] ), .IN4(n1969), .Q(
        n379) );
  AO22X1 U498 ( .IN1(n69), .IN2(n1909), .IN3(\mem[8][10] ), .IN4(n1969), .Q(
        n380) );
  AO22X1 U499 ( .IN1(n70), .IN2(n93), .IN3(\mem[8][11] ), .IN4(n1969), .Q(n381) );
  AO22X1 U500 ( .IN1(n71), .IN2(n1910), .IN3(\mem[8][12] ), .IN4(n1970), .Q(
        n382) );
  AO22X1 U501 ( .IN1(n38), .IN2(n1909), .IN3(\mem[8][13] ), .IN4(n1970), .Q(
        n383) );
  AO22X1 U502 ( .IN1(n40), .IN2(n93), .IN3(\mem[8][14] ), .IN4(n1970), .Q(n384) );
  AO22X1 U503 ( .IN1(n41), .IN2(n1910), .IN3(\mem[8][15] ), .IN4(n1970), .Q(
        n385) );
  AO22X1 U504 ( .IN1(n42), .IN2(n1909), .IN3(\mem[8][16] ), .IN4(n1970), .Q(
        n386) );
  AO22X1 U505 ( .IN1(n43), .IN2(n93), .IN3(\mem[8][17] ), .IN4(n1970), .Q(n387) );
  AO22X1 U506 ( .IN1(n44), .IN2(n1910), .IN3(\mem[8][18] ), .IN4(n1970), .Q(
        n388) );
  AO22X1 U507 ( .IN1(n45), .IN2(n1909), .IN3(\mem[8][19] ), .IN4(n1970), .Q(
        n389) );
  AO22X1 U508 ( .IN1(n46), .IN2(n93), .IN3(\mem[8][20] ), .IN4(n1970), .Q(n390) );
  AO22X1 U509 ( .IN1(n47), .IN2(n1910), .IN3(\mem[8][21] ), .IN4(n1970), .Q(
        n391) );
  AO22X1 U510 ( .IN1(n48), .IN2(n1909), .IN3(\mem[8][22] ), .IN4(n1970), .Q(
        n392) );
  AO22X1 U511 ( .IN1(n49), .IN2(n93), .IN3(\mem[8][23] ), .IN4(n1970), .Q(n393) );
  AO22X1 U512 ( .IN1(n50), .IN2(n1910), .IN3(\mem[8][24] ), .IN4(n1970), .Q(
        n394) );
  AO22X1 U513 ( .IN1(n51), .IN2(n1909), .IN3(\mem[8][25] ), .IN4(n1970), .Q(
        n395) );
  AO22X1 U514 ( .IN1(n52), .IN2(n1910), .IN3(\mem[8][26] ), .IN4(n1969), .Q(
        n396) );
  AO22X1 U515 ( .IN1(n53), .IN2(n1909), .IN3(\mem[8][27] ), .IN4(n1969), .Q(
        n397) );
  AO22X1 U516 ( .IN1(n54), .IN2(n1910), .IN3(\mem[8][28] ), .IN4(n1970), .Q(
        n398) );
  AO22X1 U517 ( .IN1(n55), .IN2(n1909), .IN3(\mem[8][29] ), .IN4(n1969), .Q(
        n399) );
  AO22X1 U518 ( .IN1(n56), .IN2(n1910), .IN3(\mem[8][30] ), .IN4(n1970), .Q(
        n400) );
  AO22X1 U519 ( .IN1(n57), .IN2(n1909), .IN3(\mem[8][31] ), .IN4(n1969), .Q(
        n401) );
  AO22X1 U521 ( .IN1(n58), .IN2(n1908), .IN3(\mem[9][0] ), .IN4(n1967), .Q(
        n402) );
  AO22X1 U522 ( .IN1(n60), .IN2(n1907), .IN3(\mem[9][1] ), .IN4(n1967), .Q(
        n403) );
  AO22X1 U523 ( .IN1(n61), .IN2(n96), .IN3(\mem[9][2] ), .IN4(n1967), .Q(n404)
         );
  AO22X1 U524 ( .IN1(n62), .IN2(n1908), .IN3(\mem[9][3] ), .IN4(n1967), .Q(
        n405) );
  AO22X1 U525 ( .IN1(n63), .IN2(n1907), .IN3(\mem[9][4] ), .IN4(n1967), .Q(
        n406) );
  AO22X1 U526 ( .IN1(n64), .IN2(n96), .IN3(\mem[9][5] ), .IN4(n1967), .Q(n407)
         );
  AO22X1 U527 ( .IN1(n65), .IN2(n1908), .IN3(\mem[9][6] ), .IN4(n1967), .Q(
        n408) );
  AO22X1 U528 ( .IN1(n66), .IN2(n1907), .IN3(\mem[9][7] ), .IN4(n1967), .Q(
        n409) );
  AO22X1 U529 ( .IN1(n67), .IN2(n96), .IN3(\mem[9][8] ), .IN4(n1967), .Q(n410)
         );
  AO22X1 U530 ( .IN1(n68), .IN2(n1908), .IN3(\mem[9][9] ), .IN4(n1967), .Q(
        n411) );
  AO22X1 U531 ( .IN1(n69), .IN2(n1907), .IN3(\mem[9][10] ), .IN4(n1967), .Q(
        n412) );
  AO22X1 U532 ( .IN1(n70), .IN2(n96), .IN3(\mem[9][11] ), .IN4(n1967), .Q(n413) );
  AO22X1 U533 ( .IN1(n71), .IN2(n1908), .IN3(\mem[9][12] ), .IN4(n1968), .Q(
        n414) );
  AO22X1 U534 ( .IN1(n1876), .IN2(n1907), .IN3(\mem[9][13] ), .IN4(n1968), .Q(
        n415) );
  AO22X1 U535 ( .IN1(n1874), .IN2(n96), .IN3(\mem[9][14] ), .IN4(n1968), .Q(
        n416) );
  AO22X1 U536 ( .IN1(n1872), .IN2(n1908), .IN3(\mem[9][15] ), .IN4(n1968), .Q(
        n417) );
  AO22X1 U537 ( .IN1(n1870), .IN2(n1907), .IN3(\mem[9][16] ), .IN4(n1968), .Q(
        n418) );
  AO22X1 U538 ( .IN1(n1868), .IN2(n96), .IN3(\mem[9][17] ), .IN4(n1968), .Q(
        n419) );
  AO22X1 U539 ( .IN1(n1866), .IN2(n1908), .IN3(\mem[9][18] ), .IN4(n1968), .Q(
        n420) );
  AO22X1 U540 ( .IN1(n1864), .IN2(n1907), .IN3(\mem[9][19] ), .IN4(n1968), .Q(
        n421) );
  AO22X1 U541 ( .IN1(n1862), .IN2(n96), .IN3(\mem[9][20] ), .IN4(n1968), .Q(
        n422) );
  AO22X1 U542 ( .IN1(n1860), .IN2(n1908), .IN3(\mem[9][21] ), .IN4(n1968), .Q(
        n423) );
  AO22X1 U543 ( .IN1(n1858), .IN2(n1907), .IN3(\mem[9][22] ), .IN4(n1968), .Q(
        n424) );
  AO22X1 U544 ( .IN1(n1856), .IN2(n96), .IN3(\mem[9][23] ), .IN4(n1968), .Q(
        n425) );
  AO22X1 U545 ( .IN1(n1854), .IN2(n1908), .IN3(\mem[9][24] ), .IN4(n1968), .Q(
        n426) );
  AO22X1 U546 ( .IN1(n1853), .IN2(n1907), .IN3(\mem[9][25] ), .IN4(n1968), .Q(
        n427) );
  AO22X1 U547 ( .IN1(n1852), .IN2(n1908), .IN3(\mem[9][26] ), .IN4(n1967), .Q(
        n428) );
  AO22X1 U548 ( .IN1(n1851), .IN2(n1907), .IN3(\mem[9][27] ), .IN4(n1968), .Q(
        n429) );
  AO22X1 U549 ( .IN1(n1850), .IN2(n1908), .IN3(\mem[9][28] ), .IN4(n1967), .Q(
        n430) );
  AO22X1 U550 ( .IN1(n1849), .IN2(n1907), .IN3(\mem[9][29] ), .IN4(n1968), .Q(
        n431) );
  AO22X1 U551 ( .IN1(n1848), .IN2(n1908), .IN3(\mem[9][30] ), .IN4(n1967), .Q(
        n432) );
  AO22X1 U552 ( .IN1(n1845), .IN2(n1907), .IN3(\mem[9][31] ), .IN4(n1967), .Q(
        n433) );
  AO22X1 U554 ( .IN1(n1844), .IN2(n1906), .IN3(\mem[10][0] ), .IN4(n1965), .Q(
        n434) );
  AO22X1 U555 ( .IN1(n1843), .IN2(n1905), .IN3(\mem[10][1] ), .IN4(n1965), .Q(
        n435) );
  AO22X1 U556 ( .IN1(n61), .IN2(n97), .IN3(\mem[10][2] ), .IN4(n1965), .Q(n436) );
  AO22X1 U557 ( .IN1(n62), .IN2(n1906), .IN3(\mem[10][3] ), .IN4(n1965), .Q(
        n437) );
  AO22X1 U558 ( .IN1(n63), .IN2(n1905), .IN3(\mem[10][4] ), .IN4(n1965), .Q(
        n438) );
  AO22X1 U559 ( .IN1(n64), .IN2(n97), .IN3(\mem[10][5] ), .IN4(n1965), .Q(n439) );
  AO22X1 U560 ( .IN1(n65), .IN2(n1906), .IN3(\mem[10][6] ), .IN4(n1965), .Q(
        n440) );
  AO22X1 U561 ( .IN1(n66), .IN2(n1905), .IN3(\mem[10][7] ), .IN4(n1965), .Q(
        n441) );
  AO22X1 U562 ( .IN1(n67), .IN2(n97), .IN3(\mem[10][8] ), .IN4(n1965), .Q(n442) );
  AO22X1 U563 ( .IN1(n68), .IN2(n1906), .IN3(\mem[10][9] ), .IN4(n1965), .Q(
        n443) );
  AO22X1 U564 ( .IN1(n69), .IN2(n1905), .IN3(\mem[10][10] ), .IN4(n1965), .Q(
        n444) );
  AO22X1 U565 ( .IN1(n70), .IN2(n97), .IN3(\mem[10][11] ), .IN4(n1965), .Q(
        n445) );
  AO22X1 U566 ( .IN1(n71), .IN2(n1906), .IN3(\mem[10][12] ), .IN4(n1966), .Q(
        n446) );
  AO22X1 U567 ( .IN1(n1875), .IN2(n1905), .IN3(\mem[10][13] ), .IN4(n1966), 
        .Q(n447) );
  AO22X1 U568 ( .IN1(n1873), .IN2(n97), .IN3(\mem[10][14] ), .IN4(n1966), .Q(
        n448) );
  AO22X1 U569 ( .IN1(n1871), .IN2(n1906), .IN3(\mem[10][15] ), .IN4(n1966), 
        .Q(n449) );
  AO22X1 U570 ( .IN1(n1869), .IN2(n1905), .IN3(\mem[10][16] ), .IN4(n1966), 
        .Q(n450) );
  AO22X1 U571 ( .IN1(n1867), .IN2(n97), .IN3(\mem[10][17] ), .IN4(n1966), .Q(
        n451) );
  AO22X1 U572 ( .IN1(n1865), .IN2(n1906), .IN3(\mem[10][18] ), .IN4(n1966), 
        .Q(n452) );
  AO22X1 U573 ( .IN1(n1863), .IN2(n1905), .IN3(\mem[10][19] ), .IN4(n1966), 
        .Q(n453) );
  AO22X1 U574 ( .IN1(n1861), .IN2(n97), .IN3(\mem[10][20] ), .IN4(n1966), .Q(
        n454) );
  AO22X1 U575 ( .IN1(n1859), .IN2(n1906), .IN3(\mem[10][21] ), .IN4(n1966), 
        .Q(n455) );
  AO22X1 U576 ( .IN1(n1857), .IN2(n1905), .IN3(\mem[10][22] ), .IN4(n1966), 
        .Q(n456) );
  AO22X1 U577 ( .IN1(n1855), .IN2(n97), .IN3(\mem[10][23] ), .IN4(n1966), .Q(
        n457) );
  AO22X1 U578 ( .IN1(n50), .IN2(n1906), .IN3(\mem[10][24] ), .IN4(n1966), .Q(
        n458) );
  AO22X1 U579 ( .IN1(n51), .IN2(n1905), .IN3(\mem[10][25] ), .IN4(n1966), .Q(
        n459) );
  AO22X1 U580 ( .IN1(n52), .IN2(n1906), .IN3(\mem[10][26] ), .IN4(n1965), .Q(
        n460) );
  AO22X1 U581 ( .IN1(n53), .IN2(n1905), .IN3(\mem[10][27] ), .IN4(n1965), .Q(
        n461) );
  AO22X1 U582 ( .IN1(n54), .IN2(n1906), .IN3(\mem[10][28] ), .IN4(n1966), .Q(
        n462) );
  AO22X1 U583 ( .IN1(n55), .IN2(n1905), .IN3(\mem[10][29] ), .IN4(n1965), .Q(
        n463) );
  AO22X1 U584 ( .IN1(n56), .IN2(n1906), .IN3(\mem[10][30] ), .IN4(n1966), .Q(
        n464) );
  AO22X1 U585 ( .IN1(n57), .IN2(n1905), .IN3(\mem[10][31] ), .IN4(n1965), .Q(
        n465) );
  AO22X1 U587 ( .IN1(n58), .IN2(n1904), .IN3(\mem[11][0] ), .IN4(n1963), .Q(
        n466) );
  AO22X1 U588 ( .IN1(n60), .IN2(n1903), .IN3(\mem[11][1] ), .IN4(n1963), .Q(
        n467) );
  AO22X1 U589 ( .IN1(n61), .IN2(n98), .IN3(\mem[11][2] ), .IN4(n1963), .Q(n468) );
  AO22X1 U590 ( .IN1(n62), .IN2(n1904), .IN3(\mem[11][3] ), .IN4(n1963), .Q(
        n469) );
  AO22X1 U591 ( .IN1(n63), .IN2(n1903), .IN3(\mem[11][4] ), .IN4(n1963), .Q(
        n470) );
  AO22X1 U592 ( .IN1(n64), .IN2(n98), .IN3(\mem[11][5] ), .IN4(n1963), .Q(n471) );
  AO22X1 U593 ( .IN1(n65), .IN2(n1904), .IN3(\mem[11][6] ), .IN4(n1963), .Q(
        n472) );
  AO22X1 U594 ( .IN1(n66), .IN2(n1903), .IN3(\mem[11][7] ), .IN4(n1963), .Q(
        n473) );
  AO22X1 U595 ( .IN1(n67), .IN2(n98), .IN3(\mem[11][8] ), .IN4(n1963), .Q(n474) );
  AO22X1 U596 ( .IN1(n68), .IN2(n1904), .IN3(\mem[11][9] ), .IN4(n1963), .Q(
        n475) );
  AO22X1 U597 ( .IN1(n69), .IN2(n1903), .IN3(\mem[11][10] ), .IN4(n1963), .Q(
        n476) );
  AO22X1 U598 ( .IN1(n70), .IN2(n98), .IN3(\mem[11][11] ), .IN4(n1963), .Q(
        n477) );
  AO22X1 U599 ( .IN1(n71), .IN2(n1904), .IN3(\mem[11][12] ), .IN4(n1964), .Q(
        n478) );
  AO22X1 U600 ( .IN1(n38), .IN2(n1903), .IN3(\mem[11][13] ), .IN4(n1964), .Q(
        n479) );
  AO22X1 U601 ( .IN1(n40), .IN2(n98), .IN3(\mem[11][14] ), .IN4(n1964), .Q(
        n480) );
  AO22X1 U602 ( .IN1(n41), .IN2(n1904), .IN3(\mem[11][15] ), .IN4(n1964), .Q(
        n481) );
  AO22X1 U603 ( .IN1(n42), .IN2(n1903), .IN3(\mem[11][16] ), .IN4(n1964), .Q(
        n482) );
  AO22X1 U604 ( .IN1(n43), .IN2(n98), .IN3(\mem[11][17] ), .IN4(n1964), .Q(
        n483) );
  AO22X1 U605 ( .IN1(n44), .IN2(n1904), .IN3(\mem[11][18] ), .IN4(n1964), .Q(
        n484) );
  AO22X1 U606 ( .IN1(n45), .IN2(n1903), .IN3(\mem[11][19] ), .IN4(n1964), .Q(
        n485) );
  AO22X1 U607 ( .IN1(n46), .IN2(n98), .IN3(\mem[11][20] ), .IN4(n1964), .Q(
        n486) );
  AO22X1 U608 ( .IN1(n47), .IN2(n1904), .IN3(\mem[11][21] ), .IN4(n1964), .Q(
        n487) );
  AO22X1 U609 ( .IN1(n48), .IN2(n1903), .IN3(\mem[11][22] ), .IN4(n1964), .Q(
        n488) );
  AO22X1 U610 ( .IN1(n49), .IN2(n98), .IN3(\mem[11][23] ), .IN4(n1964), .Q(
        n489) );
  AO22X1 U611 ( .IN1(n1854), .IN2(n1904), .IN3(\mem[11][24] ), .IN4(n1964), 
        .Q(n490) );
  AO22X1 U612 ( .IN1(n1853), .IN2(n1903), .IN3(\mem[11][25] ), .IN4(n1964), 
        .Q(n491) );
  AO22X1 U613 ( .IN1(n1852), .IN2(n1904), .IN3(\mem[11][26] ), .IN4(n1963), 
        .Q(n492) );
  AO22X1 U614 ( .IN1(n1851), .IN2(n1903), .IN3(\mem[11][27] ), .IN4(n1964), 
        .Q(n493) );
  AO22X1 U615 ( .IN1(n1850), .IN2(n1904), .IN3(\mem[11][28] ), .IN4(n1963), 
        .Q(n494) );
  AO22X1 U616 ( .IN1(n1849), .IN2(n1903), .IN3(\mem[11][29] ), .IN4(n1964), 
        .Q(n495) );
  AO22X1 U617 ( .IN1(n1848), .IN2(n1904), .IN3(\mem[11][30] ), .IN4(n1963), 
        .Q(n496) );
  AO22X1 U618 ( .IN1(n1845), .IN2(n1903), .IN3(\mem[11][31] ), .IN4(n1963), 
        .Q(n497) );
  AO22X1 U620 ( .IN1(n1844), .IN2(n1902), .IN3(\mem[12][0] ), .IN4(n1961), .Q(
        n498) );
  AO22X1 U621 ( .IN1(n1843), .IN2(n1901), .IN3(\mem[12][1] ), .IN4(n1961), .Q(
        n499) );
  AO22X1 U622 ( .IN1(n61), .IN2(n99), .IN3(\mem[12][2] ), .IN4(n1961), .Q(n500) );
  AO22X1 U623 ( .IN1(n62), .IN2(n1902), .IN3(\mem[12][3] ), .IN4(n1961), .Q(
        n501) );
  AO22X1 U624 ( .IN1(n63), .IN2(n1901), .IN3(\mem[12][4] ), .IN4(n1961), .Q(
        n502) );
  AO22X1 U625 ( .IN1(n64), .IN2(n99), .IN3(\mem[12][5] ), .IN4(n1961), .Q(n503) );
  AO22X1 U626 ( .IN1(n65), .IN2(n1902), .IN3(\mem[12][6] ), .IN4(n1961), .Q(
        n504) );
  AO22X1 U627 ( .IN1(n66), .IN2(n1901), .IN3(\mem[12][7] ), .IN4(n1961), .Q(
        n505) );
  AO22X1 U628 ( .IN1(n67), .IN2(n99), .IN3(\mem[12][8] ), .IN4(n1961), .Q(n506) );
  AO22X1 U629 ( .IN1(n68), .IN2(n1902), .IN3(\mem[12][9] ), .IN4(n1961), .Q(
        n507) );
  AO22X1 U630 ( .IN1(n69), .IN2(n1901), .IN3(\mem[12][10] ), .IN4(n1961), .Q(
        n508) );
  AO22X1 U631 ( .IN1(n70), .IN2(n99), .IN3(\mem[12][11] ), .IN4(n1961), .Q(
        n509) );
  AO22X1 U632 ( .IN1(n71), .IN2(n1902), .IN3(\mem[12][12] ), .IN4(n1962), .Q(
        n510) );
  AO22X1 U633 ( .IN1(n1876), .IN2(n1901), .IN3(\mem[12][13] ), .IN4(n1962), 
        .Q(n511) );
  AO22X1 U634 ( .IN1(n1874), .IN2(n99), .IN3(\mem[12][14] ), .IN4(n1962), .Q(
        n512) );
  AO22X1 U635 ( .IN1(n1872), .IN2(n1902), .IN3(\mem[12][15] ), .IN4(n1962), 
        .Q(n513) );
  AO22X1 U636 ( .IN1(n1870), .IN2(n1901), .IN3(\mem[12][16] ), .IN4(n1962), 
        .Q(n514) );
  AO22X1 U637 ( .IN1(n1868), .IN2(n99), .IN3(\mem[12][17] ), .IN4(n1962), .Q(
        n515) );
  AO22X1 U638 ( .IN1(n1866), .IN2(n1902), .IN3(\mem[12][18] ), .IN4(n1962), 
        .Q(n516) );
  AO22X1 U639 ( .IN1(n1864), .IN2(n1901), .IN3(\mem[12][19] ), .IN4(n1962), 
        .Q(n517) );
  AO22X1 U640 ( .IN1(n1862), .IN2(n99), .IN3(\mem[12][20] ), .IN4(n1962), .Q(
        n518) );
  AO22X1 U641 ( .IN1(n1860), .IN2(n1902), .IN3(\mem[12][21] ), .IN4(n1962), 
        .Q(n519) );
  AO22X1 U642 ( .IN1(n1858), .IN2(n1901), .IN3(\mem[12][22] ), .IN4(n1962), 
        .Q(n520) );
  AO22X1 U643 ( .IN1(n1856), .IN2(n99), .IN3(\mem[12][23] ), .IN4(n1962), .Q(
        n521) );
  AO22X1 U644 ( .IN1(n50), .IN2(n1902), .IN3(\mem[12][24] ), .IN4(n1962), .Q(
        n522) );
  AO22X1 U645 ( .IN1(n51), .IN2(n1901), .IN3(\mem[12][25] ), .IN4(n1962), .Q(
        n523) );
  AO22X1 U646 ( .IN1(n52), .IN2(n1902), .IN3(\mem[12][26] ), .IN4(n1961), .Q(
        n524) );
  AO22X1 U647 ( .IN1(n53), .IN2(n1901), .IN3(\mem[12][27] ), .IN4(n1961), .Q(
        n525) );
  AO22X1 U648 ( .IN1(n54), .IN2(n1902), .IN3(\mem[12][28] ), .IN4(n1962), .Q(
        n526) );
  AO22X1 U649 ( .IN1(n55), .IN2(n1901), .IN3(\mem[12][29] ), .IN4(n1961), .Q(
        n527) );
  AO22X1 U650 ( .IN1(n56), .IN2(n1902), .IN3(\mem[12][30] ), .IN4(n1962), .Q(
        n528) );
  AO22X1 U651 ( .IN1(n57), .IN2(n1901), .IN3(\mem[12][31] ), .IN4(n1961), .Q(
        n529) );
  AO21X1 U652 ( .IN1(n95), .IN2(n75), .IN3(n1998), .Q(n99) );
  AO22X1 U653 ( .IN1(n58), .IN2(n1900), .IN3(\mem[13][0] ), .IN4(n1959), .Q(
        n530) );
  AO22X1 U654 ( .IN1(n60), .IN2(n1899), .IN3(\mem[13][1] ), .IN4(n1959), .Q(
        n531) );
  AO22X1 U655 ( .IN1(n61), .IN2(n100), .IN3(\mem[13][2] ), .IN4(n1959), .Q(
        n532) );
  AO22X1 U656 ( .IN1(n62), .IN2(n1900), .IN3(\mem[13][3] ), .IN4(n1959), .Q(
        n533) );
  AO22X1 U657 ( .IN1(n63), .IN2(n1899), .IN3(\mem[13][4] ), .IN4(n1959), .Q(
        n534) );
  AO22X1 U658 ( .IN1(n64), .IN2(n100), .IN3(\mem[13][5] ), .IN4(n1959), .Q(
        n535) );
  AO22X1 U659 ( .IN1(n65), .IN2(n1900), .IN3(\mem[13][6] ), .IN4(n1959), .Q(
        n536) );
  AO22X1 U660 ( .IN1(n66), .IN2(n1899), .IN3(\mem[13][7] ), .IN4(n1959), .Q(
        n537) );
  AO22X1 U661 ( .IN1(n67), .IN2(n100), .IN3(\mem[13][8] ), .IN4(n1959), .Q(
        n538) );
  AO22X1 U662 ( .IN1(n68), .IN2(n1900), .IN3(\mem[13][9] ), .IN4(n1959), .Q(
        n539) );
  AO22X1 U663 ( .IN1(n69), .IN2(n1899), .IN3(\mem[13][10] ), .IN4(n1959), .Q(
        n540) );
  AO22X1 U664 ( .IN1(n70), .IN2(n100), .IN3(\mem[13][11] ), .IN4(n1959), .Q(
        n541) );
  AO22X1 U665 ( .IN1(n71), .IN2(n1900), .IN3(\mem[13][12] ), .IN4(n1960), .Q(
        n542) );
  AO22X1 U666 ( .IN1(n1875), .IN2(n1899), .IN3(\mem[13][13] ), .IN4(n1960), 
        .Q(n543) );
  AO22X1 U667 ( .IN1(n1873), .IN2(n100), .IN3(\mem[13][14] ), .IN4(n1960), .Q(
        n544) );
  AO22X1 U668 ( .IN1(n1871), .IN2(n1900), .IN3(\mem[13][15] ), .IN4(n1960), 
        .Q(n545) );
  AO22X1 U669 ( .IN1(n1869), .IN2(n1899), .IN3(\mem[13][16] ), .IN4(n1960), 
        .Q(n546) );
  AO22X1 U670 ( .IN1(n1867), .IN2(n100), .IN3(\mem[13][17] ), .IN4(n1960), .Q(
        n547) );
  AO22X1 U671 ( .IN1(n1865), .IN2(n1900), .IN3(\mem[13][18] ), .IN4(n1960), 
        .Q(n548) );
  AO22X1 U672 ( .IN1(n1863), .IN2(n1899), .IN3(\mem[13][19] ), .IN4(n1960), 
        .Q(n549) );
  AO22X1 U673 ( .IN1(n1861), .IN2(n100), .IN3(\mem[13][20] ), .IN4(n1960), .Q(
        n550) );
  AO22X1 U674 ( .IN1(n1859), .IN2(n1900), .IN3(\mem[13][21] ), .IN4(n1960), 
        .Q(n551) );
  AO22X1 U675 ( .IN1(n1857), .IN2(n1899), .IN3(\mem[13][22] ), .IN4(n1960), 
        .Q(n552) );
  AO22X1 U676 ( .IN1(n1855), .IN2(n100), .IN3(\mem[13][23] ), .IN4(n1960), .Q(
        n553) );
  AO22X1 U677 ( .IN1(n1854), .IN2(n1900), .IN3(\mem[13][24] ), .IN4(n1960), 
        .Q(n554) );
  AO22X1 U678 ( .IN1(n1853), .IN2(n1899), .IN3(\mem[13][25] ), .IN4(n1960), 
        .Q(n555) );
  AO22X1 U679 ( .IN1(n1852), .IN2(n1900), .IN3(\mem[13][26] ), .IN4(n1959), 
        .Q(n556) );
  AO22X1 U680 ( .IN1(n1851), .IN2(n1899), .IN3(\mem[13][27] ), .IN4(n1960), 
        .Q(n557) );
  AO22X1 U681 ( .IN1(n1850), .IN2(n1900), .IN3(\mem[13][28] ), .IN4(n1959), 
        .Q(n558) );
  AO22X1 U682 ( .IN1(n1849), .IN2(n1899), .IN3(\mem[13][29] ), .IN4(n1960), 
        .Q(n559) );
  AO22X1 U683 ( .IN1(n1848), .IN2(n1900), .IN3(\mem[13][30] ), .IN4(n1959), 
        .Q(n560) );
  AO22X1 U684 ( .IN1(n1845), .IN2(n1899), .IN3(\mem[13][31] ), .IN4(n1959), 
        .Q(n561) );
  AO21X1 U685 ( .IN1(n95), .IN2(n77), .IN3(n1998), .Q(n100) );
  AO22X1 U686 ( .IN1(n1844), .IN2(n1898), .IN3(\mem[14][0] ), .IN4(n1957), .Q(
        n562) );
  AO22X1 U687 ( .IN1(n1843), .IN2(n1897), .IN3(\mem[14][1] ), .IN4(n1957), .Q(
        n563) );
  AO22X1 U688 ( .IN1(n61), .IN2(n101), .IN3(\mem[14][2] ), .IN4(n1957), .Q(
        n564) );
  AO22X1 U689 ( .IN1(n62), .IN2(n1898), .IN3(\mem[14][3] ), .IN4(n1957), .Q(
        n565) );
  AO22X1 U690 ( .IN1(n63), .IN2(n1897), .IN3(\mem[14][4] ), .IN4(n1957), .Q(
        n566) );
  AO22X1 U691 ( .IN1(n64), .IN2(n101), .IN3(\mem[14][5] ), .IN4(n1957), .Q(
        n567) );
  AO22X1 U692 ( .IN1(n65), .IN2(n1898), .IN3(\mem[14][6] ), .IN4(n1957), .Q(
        n568) );
  AO22X1 U693 ( .IN1(n66), .IN2(n1897), .IN3(\mem[14][7] ), .IN4(n1957), .Q(
        n569) );
  AO22X1 U694 ( .IN1(n67), .IN2(n101), .IN3(\mem[14][8] ), .IN4(n1957), .Q(
        n570) );
  AO22X1 U695 ( .IN1(n68), .IN2(n1898), .IN3(\mem[14][9] ), .IN4(n1957), .Q(
        n571) );
  AO22X1 U696 ( .IN1(n69), .IN2(n1897), .IN3(\mem[14][10] ), .IN4(n1957), .Q(
        n572) );
  AO22X1 U697 ( .IN1(n70), .IN2(n101), .IN3(\mem[14][11] ), .IN4(n1957), .Q(
        n573) );
  AO22X1 U698 ( .IN1(n71), .IN2(n1898), .IN3(\mem[14][12] ), .IN4(n1958), .Q(
        n574) );
  AO22X1 U699 ( .IN1(n38), .IN2(n1897), .IN3(\mem[14][13] ), .IN4(n1958), .Q(
        n575) );
  AO22X1 U700 ( .IN1(n40), .IN2(n101), .IN3(\mem[14][14] ), .IN4(n1958), .Q(
        n576) );
  AO22X1 U701 ( .IN1(n41), .IN2(n1898), .IN3(\mem[14][15] ), .IN4(n1958), .Q(
        n577) );
  AO22X1 U702 ( .IN1(n42), .IN2(n1897), .IN3(\mem[14][16] ), .IN4(n1958), .Q(
        n578) );
  AO22X1 U703 ( .IN1(n43), .IN2(n101), .IN3(\mem[14][17] ), .IN4(n1958), .Q(
        n579) );
  AO22X1 U704 ( .IN1(n44), .IN2(n1898), .IN3(\mem[14][18] ), .IN4(n1958), .Q(
        n580) );
  AO22X1 U705 ( .IN1(n45), .IN2(n1897), .IN3(\mem[14][19] ), .IN4(n1958), .Q(
        n581) );
  AO22X1 U706 ( .IN1(n46), .IN2(n101), .IN3(\mem[14][20] ), .IN4(n1958), .Q(
        n582) );
  AO22X1 U707 ( .IN1(n47), .IN2(n1898), .IN3(\mem[14][21] ), .IN4(n1958), .Q(
        n583) );
  AO22X1 U708 ( .IN1(n48), .IN2(n1897), .IN3(\mem[14][22] ), .IN4(n1958), .Q(
        n584) );
  AO22X1 U709 ( .IN1(n49), .IN2(n101), .IN3(\mem[14][23] ), .IN4(n1958), .Q(
        n585) );
  AO22X1 U710 ( .IN1(n50), .IN2(n1898), .IN3(\mem[14][24] ), .IN4(n1958), .Q(
        n586) );
  AO22X1 U711 ( .IN1(n51), .IN2(n1897), .IN3(\mem[14][25] ), .IN4(n1958), .Q(
        n587) );
  AO22X1 U712 ( .IN1(n52), .IN2(n1898), .IN3(\mem[14][26] ), .IN4(n1957), .Q(
        n588) );
  AO22X1 U713 ( .IN1(n53), .IN2(n1897), .IN3(\mem[14][27] ), .IN4(n1957), .Q(
        n589) );
  AO22X1 U714 ( .IN1(n54), .IN2(n1898), .IN3(\mem[14][28] ), .IN4(n1958), .Q(
        n590) );
  AO22X1 U715 ( .IN1(n55), .IN2(n1897), .IN3(\mem[14][29] ), .IN4(n1957), .Q(
        n591) );
  AO22X1 U716 ( .IN1(n56), .IN2(n1898), .IN3(\mem[14][30] ), .IN4(n1958), .Q(
        n592) );
  AO22X1 U717 ( .IN1(n57), .IN2(n1897), .IN3(\mem[14][31] ), .IN4(n1957), .Q(
        n593) );
  AO21X1 U718 ( .IN1(n95), .IN2(n79), .IN3(n1998), .Q(n101) );
  AO22X1 U719 ( .IN1(n58), .IN2(n1896), .IN3(\mem[15][0] ), .IN4(n1955), .Q(
        n594) );
  AO22X1 U720 ( .IN1(n60), .IN2(n1895), .IN3(\mem[15][1] ), .IN4(n1955), .Q(
        n595) );
  AO22X1 U721 ( .IN1(n61), .IN2(n102), .IN3(\mem[15][2] ), .IN4(n1955), .Q(
        n596) );
  AO22X1 U722 ( .IN1(n62), .IN2(n1896), .IN3(\mem[15][3] ), .IN4(n1955), .Q(
        n597) );
  AO22X1 U723 ( .IN1(n63), .IN2(n1895), .IN3(\mem[15][4] ), .IN4(n1955), .Q(
        n598) );
  AO22X1 U724 ( .IN1(n64), .IN2(n102), .IN3(\mem[15][5] ), .IN4(n1955), .Q(
        n599) );
  AO22X1 U725 ( .IN1(n65), .IN2(n1896), .IN3(\mem[15][6] ), .IN4(n1955), .Q(
        n600) );
  AO22X1 U726 ( .IN1(n66), .IN2(n1895), .IN3(\mem[15][7] ), .IN4(n1955), .Q(
        n601) );
  AO22X1 U727 ( .IN1(n67), .IN2(n102), .IN3(\mem[15][8] ), .IN4(n1955), .Q(
        n602) );
  AO22X1 U728 ( .IN1(n68), .IN2(n1896), .IN3(\mem[15][9] ), .IN4(n1955), .Q(
        n603) );
  AO22X1 U729 ( .IN1(n69), .IN2(n1895), .IN3(\mem[15][10] ), .IN4(n1955), .Q(
        n604) );
  AO22X1 U730 ( .IN1(n70), .IN2(n102), .IN3(\mem[15][11] ), .IN4(n1955), .Q(
        n605) );
  AO22X1 U731 ( .IN1(n71), .IN2(n1896), .IN3(\mem[15][12] ), .IN4(n1956), .Q(
        n606) );
  AO22X1 U732 ( .IN1(n1876), .IN2(n1895), .IN3(\mem[15][13] ), .IN4(n1956), 
        .Q(n607) );
  AO22X1 U733 ( .IN1(n1874), .IN2(n102), .IN3(\mem[15][14] ), .IN4(n1956), .Q(
        n608) );
  AO22X1 U734 ( .IN1(n1872), .IN2(n1896), .IN3(\mem[15][15] ), .IN4(n1956), 
        .Q(n609) );
  AO22X1 U735 ( .IN1(n1870), .IN2(n1895), .IN3(\mem[15][16] ), .IN4(n1956), 
        .Q(n610) );
  AO22X1 U736 ( .IN1(n1868), .IN2(n102), .IN3(\mem[15][17] ), .IN4(n1956), .Q(
        n611) );
  AO22X1 U737 ( .IN1(n1866), .IN2(n1896), .IN3(\mem[15][18] ), .IN4(n1956), 
        .Q(n612) );
  AO22X1 U738 ( .IN1(n1864), .IN2(n1895), .IN3(\mem[15][19] ), .IN4(n1956), 
        .Q(n613) );
  AO22X1 U739 ( .IN1(n1862), .IN2(n102), .IN3(\mem[15][20] ), .IN4(n1956), .Q(
        n614) );
  AO22X1 U740 ( .IN1(n1860), .IN2(n1896), .IN3(\mem[15][21] ), .IN4(n1956), 
        .Q(n615) );
  AO22X1 U741 ( .IN1(n1858), .IN2(n1895), .IN3(\mem[15][22] ), .IN4(n1956), 
        .Q(n616) );
  AO22X1 U742 ( .IN1(n1856), .IN2(n102), .IN3(\mem[15][23] ), .IN4(n1956), .Q(
        n617) );
  AO22X1 U743 ( .IN1(n1854), .IN2(n1896), .IN3(\mem[15][24] ), .IN4(n1956), 
        .Q(n618) );
  AO22X1 U744 ( .IN1(n1853), .IN2(n1895), .IN3(\mem[15][25] ), .IN4(n1956), 
        .Q(n619) );
  AO22X1 U745 ( .IN1(n1852), .IN2(n1896), .IN3(\mem[15][26] ), .IN4(n1955), 
        .Q(n620) );
  AO22X1 U746 ( .IN1(n1851), .IN2(n1895), .IN3(\mem[15][27] ), .IN4(n1956), 
        .Q(n621) );
  AO22X1 U747 ( .IN1(n1850), .IN2(n1896), .IN3(\mem[15][28] ), .IN4(n1955), 
        .Q(n622) );
  AO22X1 U748 ( .IN1(n1849), .IN2(n1895), .IN3(\mem[15][29] ), .IN4(n1956), 
        .Q(n623) );
  AO22X1 U749 ( .IN1(n1848), .IN2(n1896), .IN3(\mem[15][30] ), .IN4(n1955), 
        .Q(n624) );
  AO22X1 U750 ( .IN1(n1845), .IN2(n1895), .IN3(\mem[15][31] ), .IN4(n1955), 
        .Q(n625) );
  AO21X1 U751 ( .IN1(n95), .IN2(n81), .IN3(n1998), .Q(n102) );
  AND3X1 U752 ( .IN1(n1836), .IN2(n2000), .IN3(wr_addr[3]), .Q(n95) );
  AO22X1 U753 ( .IN1(n1844), .IN2(n1894), .IN3(\mem[16][0] ), .IN4(n1953), .Q(
        n626) );
  AO22X1 U754 ( .IN1(n1843), .IN2(n1893), .IN3(\mem[16][1] ), .IN4(n1953), .Q(
        n627) );
  AO22X1 U755 ( .IN1(n61), .IN2(n103), .IN3(\mem[16][2] ), .IN4(n1953), .Q(
        n628) );
  AO22X1 U756 ( .IN1(n62), .IN2(n1894), .IN3(\mem[16][3] ), .IN4(n1953), .Q(
        n629) );
  AO22X1 U757 ( .IN1(n63), .IN2(n1893), .IN3(\mem[16][4] ), .IN4(n1953), .Q(
        n630) );
  AO22X1 U758 ( .IN1(n64), .IN2(n103), .IN3(\mem[16][5] ), .IN4(n1953), .Q(
        n631) );
  AO22X1 U759 ( .IN1(n65), .IN2(n1894), .IN3(\mem[16][6] ), .IN4(n1953), .Q(
        n632) );
  AO22X1 U760 ( .IN1(n66), .IN2(n1893), .IN3(\mem[16][7] ), .IN4(n1953), .Q(
        n633) );
  AO22X1 U761 ( .IN1(n67), .IN2(n103), .IN3(\mem[16][8] ), .IN4(n1953), .Q(
        n634) );
  AO22X1 U762 ( .IN1(n68), .IN2(n1894), .IN3(\mem[16][9] ), .IN4(n1953), .Q(
        n635) );
  AO22X1 U763 ( .IN1(n69), .IN2(n1893), .IN3(\mem[16][10] ), .IN4(n1953), .Q(
        n636) );
  AO22X1 U764 ( .IN1(n70), .IN2(n103), .IN3(\mem[16][11] ), .IN4(n1953), .Q(
        n637) );
  AO22X1 U765 ( .IN1(n71), .IN2(n1894), .IN3(\mem[16][12] ), .IN4(n1954), .Q(
        n638) );
  AO22X1 U766 ( .IN1(n1875), .IN2(n1893), .IN3(\mem[16][13] ), .IN4(n1954), 
        .Q(n639) );
  AO22X1 U767 ( .IN1(n1873), .IN2(n103), .IN3(\mem[16][14] ), .IN4(n1954), .Q(
        n640) );
  AO22X1 U768 ( .IN1(n1871), .IN2(n1894), .IN3(\mem[16][15] ), .IN4(n1954), 
        .Q(n641) );
  AO22X1 U769 ( .IN1(n1869), .IN2(n1893), .IN3(\mem[16][16] ), .IN4(n1954), 
        .Q(n642) );
  AO22X1 U770 ( .IN1(n1867), .IN2(n103), .IN3(\mem[16][17] ), .IN4(n1954), .Q(
        n643) );
  AO22X1 U771 ( .IN1(n1865), .IN2(n1894), .IN3(\mem[16][18] ), .IN4(n1954), 
        .Q(n644) );
  AO22X1 U772 ( .IN1(n1863), .IN2(n1893), .IN3(\mem[16][19] ), .IN4(n1954), 
        .Q(n645) );
  AO22X1 U773 ( .IN1(n1861), .IN2(n103), .IN3(\mem[16][20] ), .IN4(n1954), .Q(
        n646) );
  AO22X1 U774 ( .IN1(n1859), .IN2(n1894), .IN3(\mem[16][21] ), .IN4(n1954), 
        .Q(n647) );
  AO22X1 U775 ( .IN1(n1857), .IN2(n1893), .IN3(\mem[16][22] ), .IN4(n1954), 
        .Q(n648) );
  AO22X1 U776 ( .IN1(n1855), .IN2(n103), .IN3(\mem[16][23] ), .IN4(n1954), .Q(
        n649) );
  AO22X1 U777 ( .IN1(n50), .IN2(n1894), .IN3(\mem[16][24] ), .IN4(n1954), .Q(
        n650) );
  AO22X1 U778 ( .IN1(n51), .IN2(n1893), .IN3(\mem[16][25] ), .IN4(n1954), .Q(
        n651) );
  AO22X1 U779 ( .IN1(n52), .IN2(n1894), .IN3(\mem[16][26] ), .IN4(n1953), .Q(
        n652) );
  AO22X1 U780 ( .IN1(n53), .IN2(n1893), .IN3(\mem[16][27] ), .IN4(n1953), .Q(
        n653) );
  AO22X1 U781 ( .IN1(n54), .IN2(n1894), .IN3(\mem[16][28] ), .IN4(n1954), .Q(
        n654) );
  AO22X1 U782 ( .IN1(n55), .IN2(n1893), .IN3(\mem[16][29] ), .IN4(n1953), .Q(
        n655) );
  AO22X1 U783 ( .IN1(n56), .IN2(n1894), .IN3(\mem[16][30] ), .IN4(n1954), .Q(
        n656) );
  AO22X1 U784 ( .IN1(n57), .IN2(n1893), .IN3(\mem[16][31] ), .IN4(n1953), .Q(
        n657) );
  AO22X1 U786 ( .IN1(n58), .IN2(n1892), .IN3(\mem[17][0] ), .IN4(n1951), .Q(
        n658) );
  AO22X1 U787 ( .IN1(n60), .IN2(n1891), .IN3(\mem[17][1] ), .IN4(n1951), .Q(
        n659) );
  AO22X1 U788 ( .IN1(n61), .IN2(n105), .IN3(\mem[17][2] ), .IN4(n1951), .Q(
        n660) );
  AO22X1 U789 ( .IN1(n62), .IN2(n1892), .IN3(\mem[17][3] ), .IN4(n1951), .Q(
        n661) );
  AO22X1 U790 ( .IN1(n63), .IN2(n1891), .IN3(\mem[17][4] ), .IN4(n1951), .Q(
        n662) );
  AO22X1 U791 ( .IN1(n64), .IN2(n105), .IN3(\mem[17][5] ), .IN4(n1951), .Q(
        n663) );
  AO22X1 U792 ( .IN1(n65), .IN2(n1892), .IN3(\mem[17][6] ), .IN4(n1951), .Q(
        n664) );
  AO22X1 U793 ( .IN1(n66), .IN2(n1891), .IN3(\mem[17][7] ), .IN4(n1951), .Q(
        n665) );
  AO22X1 U794 ( .IN1(n67), .IN2(n105), .IN3(\mem[17][8] ), .IN4(n1951), .Q(
        n666) );
  AO22X1 U795 ( .IN1(n68), .IN2(n1892), .IN3(\mem[17][9] ), .IN4(n1951), .Q(
        n667) );
  AO22X1 U796 ( .IN1(n69), .IN2(n1891), .IN3(\mem[17][10] ), .IN4(n1951), .Q(
        n668) );
  AO22X1 U797 ( .IN1(n70), .IN2(n105), .IN3(\mem[17][11] ), .IN4(n1951), .Q(
        n669) );
  AO22X1 U798 ( .IN1(n71), .IN2(n1892), .IN3(\mem[17][12] ), .IN4(n1952), .Q(
        n670) );
  AO22X1 U799 ( .IN1(n38), .IN2(n1891), .IN3(\mem[17][13] ), .IN4(n1952), .Q(
        n671) );
  AO22X1 U800 ( .IN1(n40), .IN2(n105), .IN3(\mem[17][14] ), .IN4(n1952), .Q(
        n672) );
  AO22X1 U801 ( .IN1(n41), .IN2(n1892), .IN3(\mem[17][15] ), .IN4(n1952), .Q(
        n673) );
  AO22X1 U802 ( .IN1(n42), .IN2(n1891), .IN3(\mem[17][16] ), .IN4(n1952), .Q(
        n674) );
  AO22X1 U803 ( .IN1(n43), .IN2(n105), .IN3(\mem[17][17] ), .IN4(n1952), .Q(
        n675) );
  AO22X1 U804 ( .IN1(n44), .IN2(n1892), .IN3(\mem[17][18] ), .IN4(n1952), .Q(
        n676) );
  AO22X1 U805 ( .IN1(n45), .IN2(n1891), .IN3(\mem[17][19] ), .IN4(n1952), .Q(
        n677) );
  AO22X1 U806 ( .IN1(n46), .IN2(n105), .IN3(\mem[17][20] ), .IN4(n1952), .Q(
        n678) );
  AO22X1 U807 ( .IN1(n47), .IN2(n1892), .IN3(\mem[17][21] ), .IN4(n1952), .Q(
        n679) );
  AO22X1 U808 ( .IN1(n48), .IN2(n1891), .IN3(\mem[17][22] ), .IN4(n1952), .Q(
        n680) );
  AO22X1 U809 ( .IN1(n49), .IN2(n105), .IN3(\mem[17][23] ), .IN4(n1952), .Q(
        n681) );
  AO22X1 U810 ( .IN1(n1854), .IN2(n1892), .IN3(\mem[17][24] ), .IN4(n1952), 
        .Q(n682) );
  AO22X1 U811 ( .IN1(n1853), .IN2(n1891), .IN3(\mem[17][25] ), .IN4(n1952), 
        .Q(n683) );
  AO22X1 U812 ( .IN1(n1852), .IN2(n1892), .IN3(\mem[17][26] ), .IN4(n1951), 
        .Q(n684) );
  AO22X1 U813 ( .IN1(n1851), .IN2(n1891), .IN3(\mem[17][27] ), .IN4(n1952), 
        .Q(n685) );
  AO22X1 U814 ( .IN1(n1850), .IN2(n1892), .IN3(\mem[17][28] ), .IN4(n1951), 
        .Q(n686) );
  AO22X1 U815 ( .IN1(n1849), .IN2(n1891), .IN3(\mem[17][29] ), .IN4(n1952), 
        .Q(n687) );
  AO22X1 U816 ( .IN1(n1848), .IN2(n1892), .IN3(\mem[17][30] ), .IN4(n1951), 
        .Q(n688) );
  AO22X1 U817 ( .IN1(n1845), .IN2(n1891), .IN3(\mem[17][31] ), .IN4(n1951), 
        .Q(n689) );
  AO22X1 U819 ( .IN1(n1844), .IN2(n1890), .IN3(\mem[18][0] ), .IN4(n1949), .Q(
        n690) );
  AO22X1 U820 ( .IN1(n1843), .IN2(n1889), .IN3(\mem[18][1] ), .IN4(n1949), .Q(
        n691) );
  AO22X1 U821 ( .IN1(n61), .IN2(n106), .IN3(\mem[18][2] ), .IN4(n1949), .Q(
        n692) );
  AO22X1 U822 ( .IN1(n62), .IN2(n1890), .IN3(\mem[18][3] ), .IN4(n1949), .Q(
        n693) );
  AO22X1 U823 ( .IN1(n63), .IN2(n1889), .IN3(\mem[18][4] ), .IN4(n1949), .Q(
        n694) );
  AO22X1 U824 ( .IN1(n64), .IN2(n106), .IN3(\mem[18][5] ), .IN4(n1949), .Q(
        n695) );
  AO22X1 U825 ( .IN1(n65), .IN2(n1890), .IN3(\mem[18][6] ), .IN4(n1949), .Q(
        n696) );
  AO22X1 U826 ( .IN1(n66), .IN2(n1889), .IN3(\mem[18][7] ), .IN4(n1949), .Q(
        n697) );
  AO22X1 U827 ( .IN1(n67), .IN2(n106), .IN3(\mem[18][8] ), .IN4(n1949), .Q(
        n698) );
  AO22X1 U828 ( .IN1(n68), .IN2(n1890), .IN3(\mem[18][9] ), .IN4(n1949), .Q(
        n699) );
  AO22X1 U829 ( .IN1(n69), .IN2(n1889), .IN3(\mem[18][10] ), .IN4(n1949), .Q(
        n700) );
  AO22X1 U830 ( .IN1(n70), .IN2(n106), .IN3(\mem[18][11] ), .IN4(n1949), .Q(
        n701) );
  AO22X1 U831 ( .IN1(n71), .IN2(n1890), .IN3(\mem[18][12] ), .IN4(n1950), .Q(
        n702) );
  AO22X1 U832 ( .IN1(n1876), .IN2(n1889), .IN3(\mem[18][13] ), .IN4(n1950), 
        .Q(n703) );
  AO22X1 U833 ( .IN1(n1874), .IN2(n106), .IN3(\mem[18][14] ), .IN4(n1950), .Q(
        n704) );
  AO22X1 U834 ( .IN1(n1872), .IN2(n1890), .IN3(\mem[18][15] ), .IN4(n1950), 
        .Q(n705) );
  AO22X1 U835 ( .IN1(n1870), .IN2(n1889), .IN3(\mem[18][16] ), .IN4(n1950), 
        .Q(n706) );
  AO22X1 U836 ( .IN1(n1868), .IN2(n106), .IN3(\mem[18][17] ), .IN4(n1950), .Q(
        n707) );
  AO22X1 U837 ( .IN1(n1866), .IN2(n1890), .IN3(\mem[18][18] ), .IN4(n1950), 
        .Q(n708) );
  AO22X1 U838 ( .IN1(n1864), .IN2(n1889), .IN3(\mem[18][19] ), .IN4(n1950), 
        .Q(n709) );
  AO22X1 U839 ( .IN1(n1862), .IN2(n106), .IN3(\mem[18][20] ), .IN4(n1950), .Q(
        n710) );
  AO22X1 U840 ( .IN1(n1860), .IN2(n1890), .IN3(\mem[18][21] ), .IN4(n1950), 
        .Q(n711) );
  AO22X1 U841 ( .IN1(n1858), .IN2(n1889), .IN3(\mem[18][22] ), .IN4(n1950), 
        .Q(n712) );
  AO22X1 U842 ( .IN1(n1856), .IN2(n106), .IN3(\mem[18][23] ), .IN4(n1950), .Q(
        n713) );
  AO22X1 U843 ( .IN1(n50), .IN2(n1890), .IN3(\mem[18][24] ), .IN4(n1950), .Q(
        n714) );
  AO22X1 U844 ( .IN1(n51), .IN2(n1889), .IN3(\mem[18][25] ), .IN4(n1950), .Q(
        n715) );
  AO22X1 U845 ( .IN1(n52), .IN2(n1890), .IN3(\mem[18][26] ), .IN4(n1949), .Q(
        n716) );
  AO22X1 U846 ( .IN1(n53), .IN2(n1889), .IN3(\mem[18][27] ), .IN4(n1949), .Q(
        n717) );
  AO22X1 U847 ( .IN1(n54), .IN2(n1890), .IN3(\mem[18][28] ), .IN4(n1950), .Q(
        n718) );
  AO22X1 U848 ( .IN1(n55), .IN2(n1889), .IN3(\mem[18][29] ), .IN4(n1949), .Q(
        n719) );
  AO22X1 U849 ( .IN1(n56), .IN2(n1890), .IN3(\mem[18][30] ), .IN4(n1950), .Q(
        n720) );
  AO22X1 U850 ( .IN1(n57), .IN2(n1889), .IN3(\mem[18][31] ), .IN4(n1949), .Q(
        n721) );
  AO22X1 U852 ( .IN1(n58), .IN2(n1888), .IN3(\mem[19][0] ), .IN4(n1947), .Q(
        n722) );
  AO22X1 U853 ( .IN1(n60), .IN2(n1887), .IN3(\mem[19][1] ), .IN4(n1947), .Q(
        n723) );
  AO22X1 U854 ( .IN1(n61), .IN2(n107), .IN3(\mem[19][2] ), .IN4(n1947), .Q(
        n724) );
  AO22X1 U855 ( .IN1(n62), .IN2(n1888), .IN3(\mem[19][3] ), .IN4(n1947), .Q(
        n725) );
  AO22X1 U856 ( .IN1(n63), .IN2(n1887), .IN3(\mem[19][4] ), .IN4(n1947), .Q(
        n726) );
  AO22X1 U857 ( .IN1(n64), .IN2(n107), .IN3(\mem[19][5] ), .IN4(n1947), .Q(
        n727) );
  AO22X1 U858 ( .IN1(n65), .IN2(n1888), .IN3(\mem[19][6] ), .IN4(n1947), .Q(
        n728) );
  AO22X1 U859 ( .IN1(n66), .IN2(n1887), .IN3(\mem[19][7] ), .IN4(n1947), .Q(
        n729) );
  AO22X1 U860 ( .IN1(n67), .IN2(n107), .IN3(\mem[19][8] ), .IN4(n1947), .Q(
        n730) );
  AO22X1 U861 ( .IN1(n68), .IN2(n1888), .IN3(\mem[19][9] ), .IN4(n1947), .Q(
        n731) );
  AO22X1 U862 ( .IN1(n69), .IN2(n1887), .IN3(\mem[19][10] ), .IN4(n1947), .Q(
        n732) );
  AO22X1 U863 ( .IN1(n70), .IN2(n107), .IN3(\mem[19][11] ), .IN4(n1947), .Q(
        n733) );
  AO22X1 U864 ( .IN1(n71), .IN2(n1888), .IN3(\mem[19][12] ), .IN4(n1948), .Q(
        n734) );
  AO22X1 U865 ( .IN1(n1875), .IN2(n1887), .IN3(\mem[19][13] ), .IN4(n1948), 
        .Q(n735) );
  AO22X1 U866 ( .IN1(n1873), .IN2(n107), .IN3(\mem[19][14] ), .IN4(n1948), .Q(
        n736) );
  AO22X1 U867 ( .IN1(n1871), .IN2(n1888), .IN3(\mem[19][15] ), .IN4(n1948), 
        .Q(n737) );
  AO22X1 U868 ( .IN1(n1869), .IN2(n1887), .IN3(\mem[19][16] ), .IN4(n1948), 
        .Q(n738) );
  AO22X1 U869 ( .IN1(n1867), .IN2(n107), .IN3(\mem[19][17] ), .IN4(n1948), .Q(
        n739) );
  AO22X1 U870 ( .IN1(n1865), .IN2(n1888), .IN3(\mem[19][18] ), .IN4(n1948), 
        .Q(n740) );
  AO22X1 U871 ( .IN1(n1863), .IN2(n1887), .IN3(\mem[19][19] ), .IN4(n1948), 
        .Q(n741) );
  AO22X1 U872 ( .IN1(n1861), .IN2(n107), .IN3(\mem[19][20] ), .IN4(n1948), .Q(
        n742) );
  AO22X1 U873 ( .IN1(n1859), .IN2(n1888), .IN3(\mem[19][21] ), .IN4(n1948), 
        .Q(n743) );
  AO22X1 U874 ( .IN1(n1857), .IN2(n1887), .IN3(\mem[19][22] ), .IN4(n1948), 
        .Q(n744) );
  AO22X1 U875 ( .IN1(n1855), .IN2(n107), .IN3(\mem[19][23] ), .IN4(n1948), .Q(
        n745) );
  AO22X1 U876 ( .IN1(n1854), .IN2(n1888), .IN3(\mem[19][24] ), .IN4(n1948), 
        .Q(n746) );
  AO22X1 U877 ( .IN1(n1853), .IN2(n1887), .IN3(\mem[19][25] ), .IN4(n1948), 
        .Q(n747) );
  AO22X1 U878 ( .IN1(n1852), .IN2(n1888), .IN3(\mem[19][26] ), .IN4(n1947), 
        .Q(n748) );
  AO22X1 U879 ( .IN1(n1851), .IN2(n1887), .IN3(\mem[19][27] ), .IN4(n1948), 
        .Q(n749) );
  AO22X1 U880 ( .IN1(n1850), .IN2(n1888), .IN3(\mem[19][28] ), .IN4(n1947), 
        .Q(n750) );
  AO22X1 U881 ( .IN1(n1849), .IN2(n1887), .IN3(\mem[19][29] ), .IN4(n1948), 
        .Q(n751) );
  AO22X1 U882 ( .IN1(n1848), .IN2(n1888), .IN3(\mem[19][30] ), .IN4(n1947), 
        .Q(n752) );
  AO22X1 U883 ( .IN1(n1845), .IN2(n1887), .IN3(\mem[19][31] ), .IN4(n1947), 
        .Q(n753) );
  AND3X1 U885 ( .IN1(wr_addr[1]), .IN2(n2002), .IN3(wr_addr[0]), .Q(n72) );
  AO22X1 U886 ( .IN1(n1844), .IN2(n1886), .IN3(\mem[20][0] ), .IN4(n1945), .Q(
        n754) );
  AO22X1 U887 ( .IN1(n1843), .IN2(n1885), .IN3(\mem[20][1] ), .IN4(n1945), .Q(
        n755) );
  AO22X1 U888 ( .IN1(n61), .IN2(n108), .IN3(\mem[20][2] ), .IN4(n1945), .Q(
        n756) );
  AO22X1 U889 ( .IN1(n62), .IN2(n1886), .IN3(\mem[20][3] ), .IN4(n1945), .Q(
        n757) );
  AO22X1 U890 ( .IN1(n63), .IN2(n1885), .IN3(\mem[20][4] ), .IN4(n1945), .Q(
        n758) );
  AO22X1 U891 ( .IN1(n64), .IN2(n108), .IN3(\mem[20][5] ), .IN4(n1945), .Q(
        n759) );
  AO22X1 U892 ( .IN1(n65), .IN2(n1886), .IN3(\mem[20][6] ), .IN4(n1945), .Q(
        n760) );
  AO22X1 U893 ( .IN1(n66), .IN2(n1885), .IN3(\mem[20][7] ), .IN4(n1945), .Q(
        n761) );
  AO22X1 U894 ( .IN1(n67), .IN2(n108), .IN3(\mem[20][8] ), .IN4(n1945), .Q(
        n762) );
  AO22X1 U895 ( .IN1(n68), .IN2(n1886), .IN3(\mem[20][9] ), .IN4(n1945), .Q(
        n763) );
  AO22X1 U896 ( .IN1(n69), .IN2(n1885), .IN3(\mem[20][10] ), .IN4(n1945), .Q(
        n764) );
  AO22X1 U897 ( .IN1(n70), .IN2(n108), .IN3(\mem[20][11] ), .IN4(n1945), .Q(
        n765) );
  AO22X1 U898 ( .IN1(n71), .IN2(n1886), .IN3(\mem[20][12] ), .IN4(n1946), .Q(
        n766) );
  AO22X1 U899 ( .IN1(n38), .IN2(n1885), .IN3(\mem[20][13] ), .IN4(n1946), .Q(
        n767) );
  AO22X1 U900 ( .IN1(n40), .IN2(n108), .IN3(\mem[20][14] ), .IN4(n1946), .Q(
        n768) );
  AO22X1 U901 ( .IN1(n41), .IN2(n1886), .IN3(\mem[20][15] ), .IN4(n1946), .Q(
        n769) );
  AO22X1 U902 ( .IN1(n42), .IN2(n1885), .IN3(\mem[20][16] ), .IN4(n1946), .Q(
        n770) );
  AO22X1 U903 ( .IN1(n43), .IN2(n108), .IN3(\mem[20][17] ), .IN4(n1946), .Q(
        n771) );
  AO22X1 U904 ( .IN1(n44), .IN2(n1886), .IN3(\mem[20][18] ), .IN4(n1946), .Q(
        n772) );
  AO22X1 U905 ( .IN1(n45), .IN2(n1885), .IN3(\mem[20][19] ), .IN4(n1946), .Q(
        n773) );
  AO22X1 U906 ( .IN1(n46), .IN2(n108), .IN3(\mem[20][20] ), .IN4(n1946), .Q(
        n774) );
  AO22X1 U907 ( .IN1(n47), .IN2(n1886), .IN3(\mem[20][21] ), .IN4(n1946), .Q(
        n775) );
  AO22X1 U908 ( .IN1(n48), .IN2(n1885), .IN3(\mem[20][22] ), .IN4(n1946), .Q(
        n776) );
  AO22X1 U909 ( .IN1(n49), .IN2(n108), .IN3(\mem[20][23] ), .IN4(n1946), .Q(
        n777) );
  AO22X1 U910 ( .IN1(n50), .IN2(n1886), .IN3(\mem[20][24] ), .IN4(n1946), .Q(
        n778) );
  AO22X1 U911 ( .IN1(n51), .IN2(n1885), .IN3(\mem[20][25] ), .IN4(n1946), .Q(
        n779) );
  AO22X1 U912 ( .IN1(n52), .IN2(n1886), .IN3(\mem[20][26] ), .IN4(n1945), .Q(
        n780) );
  AO22X1 U913 ( .IN1(n53), .IN2(n1885), .IN3(\mem[20][27] ), .IN4(n1945), .Q(
        n781) );
  AO22X1 U914 ( .IN1(n54), .IN2(n1886), .IN3(\mem[20][28] ), .IN4(n1946), .Q(
        n782) );
  AO22X1 U915 ( .IN1(n55), .IN2(n1885), .IN3(\mem[20][29] ), .IN4(n1945), .Q(
        n783) );
  AO22X1 U916 ( .IN1(n56), .IN2(n1886), .IN3(\mem[20][30] ), .IN4(n1946), .Q(
        n784) );
  AO22X1 U917 ( .IN1(n57), .IN2(n1885), .IN3(\mem[20][31] ), .IN4(n1945), .Q(
        n785) );
  AO21X1 U918 ( .IN1(n104), .IN2(n75), .IN3(n1999), .Q(n108) );
  AND3X1 U919 ( .IN1(n2004), .IN2(n2003), .IN3(wr_addr[2]), .Q(n75) );
  AO22X1 U920 ( .IN1(n58), .IN2(n1884), .IN3(\mem[21][0] ), .IN4(n1943), .Q(
        n786) );
  AO22X1 U921 ( .IN1(n60), .IN2(n1883), .IN3(\mem[21][1] ), .IN4(n1943), .Q(
        n787) );
  AO22X1 U922 ( .IN1(n61), .IN2(n109), .IN3(\mem[21][2] ), .IN4(n1943), .Q(
        n788) );
  AO22X1 U923 ( .IN1(n62), .IN2(n1884), .IN3(\mem[21][3] ), .IN4(n1943), .Q(
        n789) );
  AO22X1 U924 ( .IN1(n63), .IN2(n1883), .IN3(\mem[21][4] ), .IN4(n1943), .Q(
        n790) );
  AO22X1 U925 ( .IN1(n64), .IN2(n109), .IN3(\mem[21][5] ), .IN4(n1943), .Q(
        n791) );
  AO22X1 U926 ( .IN1(n65), .IN2(n1884), .IN3(\mem[21][6] ), .IN4(n1943), .Q(
        n792) );
  AO22X1 U927 ( .IN1(n66), .IN2(n1883), .IN3(\mem[21][7] ), .IN4(n1943), .Q(
        n793) );
  AO22X1 U928 ( .IN1(n67), .IN2(n109), .IN3(\mem[21][8] ), .IN4(n1943), .Q(
        n794) );
  AO22X1 U929 ( .IN1(n68), .IN2(n1884), .IN3(\mem[21][9] ), .IN4(n1943), .Q(
        n795) );
  AO22X1 U930 ( .IN1(n69), .IN2(n1883), .IN3(\mem[21][10] ), .IN4(n1943), .Q(
        n796) );
  AO22X1 U931 ( .IN1(n70), .IN2(n109), .IN3(\mem[21][11] ), .IN4(n1943), .Q(
        n797) );
  AO22X1 U932 ( .IN1(n71), .IN2(n1884), .IN3(\mem[21][12] ), .IN4(n1944), .Q(
        n798) );
  AO22X1 U933 ( .IN1(n1876), .IN2(n1883), .IN3(\mem[21][13] ), .IN4(n1944), 
        .Q(n799) );
  AO22X1 U934 ( .IN1(n1874), .IN2(n109), .IN3(\mem[21][14] ), .IN4(n1944), .Q(
        n800) );
  AO22X1 U935 ( .IN1(n1872), .IN2(n1884), .IN3(\mem[21][15] ), .IN4(n1944), 
        .Q(n801) );
  AO22X1 U936 ( .IN1(n1870), .IN2(n1883), .IN3(\mem[21][16] ), .IN4(n1944), 
        .Q(n802) );
  AO22X1 U937 ( .IN1(n1868), .IN2(n109), .IN3(\mem[21][17] ), .IN4(n1944), .Q(
        n803) );
  AO22X1 U938 ( .IN1(n1866), .IN2(n1884), .IN3(\mem[21][18] ), .IN4(n1944), 
        .Q(n804) );
  AO22X1 U939 ( .IN1(n1864), .IN2(n1883), .IN3(\mem[21][19] ), .IN4(n1944), 
        .Q(n805) );
  AO22X1 U940 ( .IN1(n1862), .IN2(n109), .IN3(\mem[21][20] ), .IN4(n1944), .Q(
        n806) );
  AO22X1 U941 ( .IN1(n1860), .IN2(n1884), .IN3(\mem[21][21] ), .IN4(n1944), 
        .Q(n807) );
  AO22X1 U942 ( .IN1(n1858), .IN2(n1883), .IN3(\mem[21][22] ), .IN4(n1944), 
        .Q(n808) );
  AO22X1 U943 ( .IN1(n1856), .IN2(n109), .IN3(\mem[21][23] ), .IN4(n1944), .Q(
        n809) );
  AO22X1 U944 ( .IN1(n1854), .IN2(n1884), .IN3(\mem[21][24] ), .IN4(n1944), 
        .Q(n810) );
  AO22X1 U945 ( .IN1(n1853), .IN2(n1883), .IN3(\mem[21][25] ), .IN4(n1944), 
        .Q(n811) );
  AO22X1 U946 ( .IN1(n1852), .IN2(n1884), .IN3(\mem[21][26] ), .IN4(n1943), 
        .Q(n812) );
  AO22X1 U947 ( .IN1(n1851), .IN2(n1883), .IN3(\mem[21][27] ), .IN4(n1944), 
        .Q(n813) );
  AO22X1 U948 ( .IN1(n1850), .IN2(n1884), .IN3(\mem[21][28] ), .IN4(n1943), 
        .Q(n814) );
  AO22X1 U949 ( .IN1(n1849), .IN2(n1883), .IN3(\mem[21][29] ), .IN4(n1944), 
        .Q(n815) );
  AO22X1 U950 ( .IN1(n1848), .IN2(n1884), .IN3(\mem[21][30] ), .IN4(n1943), 
        .Q(n816) );
  AO22X1 U951 ( .IN1(n1845), .IN2(n1883), .IN3(\mem[21][31] ), .IN4(n1943), 
        .Q(n817) );
  AO21X1 U952 ( .IN1(n104), .IN2(n77), .IN3(n1999), .Q(n109) );
  AND3X1 U953 ( .IN1(wr_addr[0]), .IN2(n2003), .IN3(wr_addr[2]), .Q(n77) );
  AO22X1 U954 ( .IN1(n1844), .IN2(n1882), .IN3(\mem[22][0] ), .IN4(n1941), .Q(
        n818) );
  AO22X1 U955 ( .IN1(n1843), .IN2(n1881), .IN3(\mem[22][1] ), .IN4(n1941), .Q(
        n819) );
  AO22X1 U956 ( .IN1(n61), .IN2(n110), .IN3(\mem[22][2] ), .IN4(n1941), .Q(
        n820) );
  AO22X1 U957 ( .IN1(n62), .IN2(n1882), .IN3(\mem[22][3] ), .IN4(n1941), .Q(
        n821) );
  AO22X1 U958 ( .IN1(n63), .IN2(n1881), .IN3(\mem[22][4] ), .IN4(n1941), .Q(
        n822) );
  AO22X1 U959 ( .IN1(n64), .IN2(n110), .IN3(\mem[22][5] ), .IN4(n1941), .Q(
        n823) );
  AO22X1 U960 ( .IN1(n65), .IN2(n1882), .IN3(\mem[22][6] ), .IN4(n1941), .Q(
        n824) );
  AO22X1 U961 ( .IN1(n66), .IN2(n1881), .IN3(\mem[22][7] ), .IN4(n1941), .Q(
        n825) );
  AO22X1 U962 ( .IN1(n67), .IN2(n110), .IN3(\mem[22][8] ), .IN4(n1941), .Q(
        n826) );
  AO22X1 U963 ( .IN1(n68), .IN2(n1882), .IN3(\mem[22][9] ), .IN4(n1941), .Q(
        n827) );
  AO22X1 U964 ( .IN1(n69), .IN2(n1881), .IN3(\mem[22][10] ), .IN4(n1941), .Q(
        n828) );
  AO22X1 U965 ( .IN1(n70), .IN2(n110), .IN3(\mem[22][11] ), .IN4(n1941), .Q(
        n829) );
  AO22X1 U966 ( .IN1(n71), .IN2(n1882), .IN3(\mem[22][12] ), .IN4(n1942), .Q(
        n830) );
  AO22X1 U967 ( .IN1(n1875), .IN2(n1881), .IN3(\mem[22][13] ), .IN4(n1942), 
        .Q(n831) );
  AO22X1 U968 ( .IN1(n1873), .IN2(n110), .IN3(\mem[22][14] ), .IN4(n1942), .Q(
        n832) );
  AO22X1 U969 ( .IN1(n1871), .IN2(n1882), .IN3(\mem[22][15] ), .IN4(n1942), 
        .Q(n833) );
  AO22X1 U970 ( .IN1(n1869), .IN2(n1881), .IN3(\mem[22][16] ), .IN4(n1942), 
        .Q(n834) );
  AO22X1 U971 ( .IN1(n1867), .IN2(n110), .IN3(\mem[22][17] ), .IN4(n1942), .Q(
        n835) );
  AO22X1 U972 ( .IN1(n1865), .IN2(n1882), .IN3(\mem[22][18] ), .IN4(n1942), 
        .Q(n836) );
  AO22X1 U973 ( .IN1(n1863), .IN2(n1881), .IN3(\mem[22][19] ), .IN4(n1942), 
        .Q(n837) );
  AO22X1 U974 ( .IN1(n1861), .IN2(n110), .IN3(\mem[22][20] ), .IN4(n1942), .Q(
        n838) );
  AO22X1 U975 ( .IN1(n1859), .IN2(n1882), .IN3(\mem[22][21] ), .IN4(n1942), 
        .Q(n839) );
  AO22X1 U976 ( .IN1(n1857), .IN2(n1881), .IN3(\mem[22][22] ), .IN4(n1942), 
        .Q(n840) );
  AO22X1 U977 ( .IN1(n1855), .IN2(n110), .IN3(\mem[22][23] ), .IN4(n1942), .Q(
        n841) );
  AO22X1 U978 ( .IN1(n50), .IN2(n1882), .IN3(\mem[22][24] ), .IN4(n1942), .Q(
        n842) );
  AO22X1 U979 ( .IN1(n51), .IN2(n1881), .IN3(\mem[22][25] ), .IN4(n1942), .Q(
        n843) );
  AO22X1 U980 ( .IN1(n52), .IN2(n1882), .IN3(\mem[22][26] ), .IN4(n1941), .Q(
        n844) );
  AO22X1 U981 ( .IN1(n53), .IN2(n1881), .IN3(\mem[22][27] ), .IN4(n1941), .Q(
        n845) );
  AO22X1 U982 ( .IN1(n54), .IN2(n1882), .IN3(\mem[22][28] ), .IN4(n1942), .Q(
        n846) );
  AO22X1 U983 ( .IN1(n55), .IN2(n1881), .IN3(\mem[22][29] ), .IN4(n1941), .Q(
        n847) );
  AO22X1 U984 ( .IN1(n56), .IN2(n1882), .IN3(\mem[22][30] ), .IN4(n1942), .Q(
        n848) );
  AO22X1 U985 ( .IN1(n57), .IN2(n1881), .IN3(\mem[22][31] ), .IN4(n1941), .Q(
        n849) );
  AO21X1 U986 ( .IN1(n104), .IN2(n79), .IN3(n1999), .Q(n110) );
  AND3X1 U987 ( .IN1(wr_addr[1]), .IN2(n2004), .IN3(wr_addr[2]), .Q(n79) );
  AO22X1 U988 ( .IN1(n58), .IN2(n1880), .IN3(\mem[23][0] ), .IN4(n1939), .Q(
        n850) );
  AO22X1 U989 ( .IN1(n60), .IN2(n1879), .IN3(\mem[23][1] ), .IN4(n1939), .Q(
        n851) );
  AO22X1 U990 ( .IN1(n61), .IN2(n111), .IN3(\mem[23][2] ), .IN4(n1939), .Q(
        n852) );
  AO22X1 U991 ( .IN1(n62), .IN2(n1880), .IN3(\mem[23][3] ), .IN4(n1939), .Q(
        n853) );
  AO22X1 U992 ( .IN1(n63), .IN2(n1879), .IN3(\mem[23][4] ), .IN4(n1939), .Q(
        n854) );
  AO22X1 U993 ( .IN1(n64), .IN2(n111), .IN3(\mem[23][5] ), .IN4(n1939), .Q(
        n855) );
  AO22X1 U994 ( .IN1(n65), .IN2(n1880), .IN3(\mem[23][6] ), .IN4(n1939), .Q(
        n856) );
  AO22X1 U995 ( .IN1(n66), .IN2(n1879), .IN3(\mem[23][7] ), .IN4(n1939), .Q(
        n857) );
  AO22X1 U996 ( .IN1(n67), .IN2(n111), .IN3(\mem[23][8] ), .IN4(n1939), .Q(
        n858) );
  AO22X1 U997 ( .IN1(n68), .IN2(n1880), .IN3(\mem[23][9] ), .IN4(n1939), .Q(
        n859) );
  AO22X1 U998 ( .IN1(n69), .IN2(n1879), .IN3(\mem[23][10] ), .IN4(n1939), .Q(
        n860) );
  AO22X1 U999 ( .IN1(n70), .IN2(n111), .IN3(\mem[23][11] ), .IN4(n1939), .Q(
        n861) );
  AO22X1 U1000 ( .IN1(n71), .IN2(n1880), .IN3(\mem[23][12] ), .IN4(n1940), .Q(
        n862) );
  AO22X1 U1001 ( .IN1(n38), .IN2(n1879), .IN3(\mem[23][13] ), .IN4(n1940), .Q(
        n863) );
  AO22X1 U1002 ( .IN1(n40), .IN2(n111), .IN3(\mem[23][14] ), .IN4(n1940), .Q(
        n864) );
  AO22X1 U1003 ( .IN1(n41), .IN2(n1880), .IN3(\mem[23][15] ), .IN4(n1940), .Q(
        n865) );
  AO22X1 U1004 ( .IN1(n42), .IN2(n1879), .IN3(\mem[23][16] ), .IN4(n1940), .Q(
        n866) );
  AO22X1 U1005 ( .IN1(n43), .IN2(n111), .IN3(\mem[23][17] ), .IN4(n1940), .Q(
        n867) );
  AO22X1 U1006 ( .IN1(n44), .IN2(n1880), .IN3(\mem[23][18] ), .IN4(n1940), .Q(
        n868) );
  AO22X1 U1007 ( .IN1(n45), .IN2(n1879), .IN3(\mem[23][19] ), .IN4(n1940), .Q(
        n869) );
  AO22X1 U1008 ( .IN1(n46), .IN2(n111), .IN3(\mem[23][20] ), .IN4(n1940), .Q(
        n870) );
  AO22X1 U1009 ( .IN1(n47), .IN2(n1880), .IN3(\mem[23][21] ), .IN4(n1940), .Q(
        n871) );
  AO22X1 U1010 ( .IN1(n48), .IN2(n1879), .IN3(\mem[23][22] ), .IN4(n1940), .Q(
        n872) );
  AO22X1 U1011 ( .IN1(n49), .IN2(n111), .IN3(\mem[23][23] ), .IN4(n1940), .Q(
        n873) );
  AO22X1 U1012 ( .IN1(n1854), .IN2(n1880), .IN3(\mem[23][24] ), .IN4(n1940), 
        .Q(n874) );
  AO22X1 U1013 ( .IN1(n1853), .IN2(n1879), .IN3(\mem[23][25] ), .IN4(n1940), 
        .Q(n875) );
  AO22X1 U1014 ( .IN1(n1852), .IN2(n1880), .IN3(\mem[23][26] ), .IN4(n1939), 
        .Q(n876) );
  AO22X1 U1015 ( .IN1(n1851), .IN2(n1879), .IN3(\mem[23][27] ), .IN4(n1940), 
        .Q(n877) );
  AO22X1 U1016 ( .IN1(n1850), .IN2(n1880), .IN3(\mem[23][28] ), .IN4(n1939), 
        .Q(n878) );
  AO22X1 U1017 ( .IN1(n1849), .IN2(n1879), .IN3(\mem[23][29] ), .IN4(n1940), 
        .Q(n879) );
  AO22X1 U1018 ( .IN1(n1848), .IN2(n1880), .IN3(\mem[23][30] ), .IN4(n1939), 
        .Q(n880) );
  AO22X1 U1019 ( .IN1(n1845), .IN2(n1879), .IN3(\mem[23][31] ), .IN4(n1939), 
        .Q(n881) );
  AO21X1 U1020 ( .IN1(n104), .IN2(n81), .IN3(n1999), .Q(n111) );
  AND3X1 U1021 ( .IN1(wr_addr[0]), .IN2(wr_addr[1]), .IN3(wr_addr[2]), .Q(n81)
         );
  AND3X1 U1022 ( .IN1(n1835), .IN2(n2001), .IN3(wr_addr[4]), .Q(n104) );
  AO22X1 U1023 ( .IN1(n1844), .IN2(n1878), .IN3(\mem[24][0] ), .IN4(n1937), 
        .Q(n882) );
  AO22X1 U1024 ( .IN1(n1843), .IN2(n1877), .IN3(\mem[24][1] ), .IN4(n1937), 
        .Q(n883) );
  AO22X1 U1025 ( .IN1(n61), .IN2(n112), .IN3(\mem[24][2] ), .IN4(n1937), .Q(
        n884) );
  AO22X1 U1026 ( .IN1(n62), .IN2(n1878), .IN3(\mem[24][3] ), .IN4(n1937), .Q(
        n885) );
  AO22X1 U1027 ( .IN1(n63), .IN2(n1877), .IN3(\mem[24][4] ), .IN4(n1937), .Q(
        n886) );
  AO22X1 U1028 ( .IN1(n64), .IN2(n112), .IN3(\mem[24][5] ), .IN4(n1937), .Q(
        n887) );
  AO22X1 U1029 ( .IN1(n65), .IN2(n1878), .IN3(\mem[24][6] ), .IN4(n1937), .Q(
        n888) );
  AO22X1 U1030 ( .IN1(n66), .IN2(n1877), .IN3(\mem[24][7] ), .IN4(n1937), .Q(
        n889) );
  AO22X1 U1031 ( .IN1(n67), .IN2(n112), .IN3(\mem[24][8] ), .IN4(n1937), .Q(
        n890) );
  AO22X1 U1032 ( .IN1(n68), .IN2(n1878), .IN3(\mem[24][9] ), .IN4(n1937), .Q(
        n891) );
  AO22X1 U1033 ( .IN1(n69), .IN2(n1877), .IN3(\mem[24][10] ), .IN4(n1937), .Q(
        n892) );
  AO22X1 U1034 ( .IN1(n70), .IN2(n112), .IN3(\mem[24][11] ), .IN4(n1937), .Q(
        n893) );
  AO22X1 U1035 ( .IN1(n71), .IN2(n1878), .IN3(\mem[24][12] ), .IN4(n1938), .Q(
        n894) );
  AO22X1 U1036 ( .IN1(n1876), .IN2(n1877), .IN3(\mem[24][13] ), .IN4(n1938), 
        .Q(n895) );
  AO22X1 U1037 ( .IN1(n1874), .IN2(n112), .IN3(\mem[24][14] ), .IN4(n1938), 
        .Q(n896) );
  AO22X1 U1038 ( .IN1(n1872), .IN2(n1878), .IN3(\mem[24][15] ), .IN4(n1938), 
        .Q(n897) );
  AO22X1 U1039 ( .IN1(n1870), .IN2(n1877), .IN3(\mem[24][16] ), .IN4(n1938), 
        .Q(n898) );
  AO22X1 U1040 ( .IN1(n1868), .IN2(n112), .IN3(\mem[24][17] ), .IN4(n1938), 
        .Q(n899) );
  AO22X1 U1041 ( .IN1(n1866), .IN2(n1878), .IN3(\mem[24][18] ), .IN4(n1938), 
        .Q(n900) );
  AO22X1 U1042 ( .IN1(n1864), .IN2(n1877), .IN3(\mem[24][19] ), .IN4(n1938), 
        .Q(n901) );
  AO22X1 U1043 ( .IN1(n1862), .IN2(n112), .IN3(\mem[24][20] ), .IN4(n1938), 
        .Q(n902) );
  AO22X1 U1044 ( .IN1(n1860), .IN2(n1878), .IN3(\mem[24][21] ), .IN4(n1938), 
        .Q(n903) );
  AO22X1 U1045 ( .IN1(n1858), .IN2(n1877), .IN3(\mem[24][22] ), .IN4(n1938), 
        .Q(n904) );
  AO22X1 U1046 ( .IN1(n1856), .IN2(n112), .IN3(\mem[24][23] ), .IN4(n1938), 
        .Q(n905) );
  AO22X1 U1047 ( .IN1(n50), .IN2(n1878), .IN3(\mem[24][24] ), .IN4(n1938), .Q(
        n906) );
  AO22X1 U1048 ( .IN1(n51), .IN2(n1877), .IN3(\mem[24][25] ), .IN4(n1938), .Q(
        n907) );
  AO22X1 U1049 ( .IN1(n52), .IN2(n1878), .IN3(\mem[24][26] ), .IN4(n1937), .Q(
        n908) );
  AO22X1 U1050 ( .IN1(n53), .IN2(n1877), .IN3(\mem[24][27] ), .IN4(n1937), .Q(
        n909) );
  AO22X1 U1051 ( .IN1(n54), .IN2(n1878), .IN3(\mem[24][28] ), .IN4(n1938), .Q(
        n910) );
  AO22X1 U1052 ( .IN1(n55), .IN2(n1877), .IN3(\mem[24][29] ), .IN4(n1937), .Q(
        n911) );
  AO22X1 U1053 ( .IN1(n56), .IN2(n1878), .IN3(\mem[24][30] ), .IN4(n1938), .Q(
        n912) );
  AO22X1 U1054 ( .IN1(n57), .IN2(n1877), .IN3(\mem[24][31] ), .IN4(n1937), .Q(
        n913) );
  AO21X1 U1055 ( .IN1(n94), .IN2(n73), .IN3(n1999), .Q(n112) );
  AND3X1 U1056 ( .IN1(n2003), .IN2(n2002), .IN3(n2004), .Q(n94) );
  AO22X1 U1057 ( .IN1(n58), .IN2(n1847), .IN3(\mem[25][0] ), .IN4(n1935), .Q(
        n914) );
  AO22X1 U1058 ( .IN1(n60), .IN2(n1846), .IN3(\mem[25][1] ), .IN4(n1935), .Q(
        n915) );
  AO22X1 U1059 ( .IN1(n61), .IN2(n113), .IN3(\mem[25][2] ), .IN4(n1935), .Q(
        n916) );
  AO22X1 U1060 ( .IN1(n62), .IN2(n1847), .IN3(\mem[25][3] ), .IN4(n1935), .Q(
        n917) );
  AO22X1 U1061 ( .IN1(n63), .IN2(n1846), .IN3(\mem[25][4] ), .IN4(n1935), .Q(
        n918) );
  AO22X1 U1062 ( .IN1(n64), .IN2(n113), .IN3(\mem[25][5] ), .IN4(n1935), .Q(
        n919) );
  AO22X1 U1063 ( .IN1(n65), .IN2(n1847), .IN3(\mem[25][6] ), .IN4(n1935), .Q(
        n920) );
  AO22X1 U1064 ( .IN1(n66), .IN2(n1846), .IN3(\mem[25][7] ), .IN4(n1935), .Q(
        n921) );
  AO22X1 U1065 ( .IN1(n67), .IN2(n113), .IN3(\mem[25][8] ), .IN4(n1935), .Q(
        n922) );
  AO22X1 U1066 ( .IN1(n68), .IN2(n1847), .IN3(\mem[25][9] ), .IN4(n1935), .Q(
        n923) );
  AO22X1 U1067 ( .IN1(n69), .IN2(n1846), .IN3(\mem[25][10] ), .IN4(n1935), .Q(
        n924) );
  AO22X1 U1068 ( .IN1(n70), .IN2(n113), .IN3(\mem[25][11] ), .IN4(n1935), .Q(
        n925) );
  AO22X1 U1069 ( .IN1(n71), .IN2(n1847), .IN3(\mem[25][12] ), .IN4(n1936), .Q(
        n926) );
  AO22X1 U1070 ( .IN1(n1875), .IN2(n1846), .IN3(\mem[25][13] ), .IN4(n1936), 
        .Q(n927) );
  AO22X1 U1072 ( .IN1(n1873), .IN2(n113), .IN3(\mem[25][14] ), .IN4(n1936), 
        .Q(n928) );
  AO22X1 U1074 ( .IN1(n1871), .IN2(n1847), .IN3(\mem[25][15] ), .IN4(n1936), 
        .Q(n929) );
  AO22X1 U1076 ( .IN1(n1869), .IN2(n1846), .IN3(\mem[25][16] ), .IN4(n1936), 
        .Q(n930) );
  AND2X1 U1077 ( .IN1(wr_data[16]), .IN2(n1836), .Q(n42) );
  AO22X1 U1078 ( .IN1(n1867), .IN2(n113), .IN3(\mem[25][17] ), .IN4(n1936), 
        .Q(n931) );
  AND2X1 U1079 ( .IN1(wr_data[17]), .IN2(n1835), .Q(n43) );
  AO22X1 U1080 ( .IN1(n1865), .IN2(n1847), .IN3(\mem[25][18] ), .IN4(n1936), 
        .Q(n932) );
  AND2X1 U1081 ( .IN1(wr_data[18]), .IN2(n1836), .Q(n44) );
  AO22X1 U1082 ( .IN1(n1863), .IN2(n1846), .IN3(\mem[25][19] ), .IN4(n1936), 
        .Q(n933) );
  AND2X1 U1083 ( .IN1(wr_data[19]), .IN2(n1835), .Q(n45) );
  AO22X1 U1084 ( .IN1(n1861), .IN2(n113), .IN3(\mem[25][20] ), .IN4(n1936), 
        .Q(n934) );
  AND2X1 U1085 ( .IN1(wr_data[20]), .IN2(n1838), .Q(n46) );
  AO22X1 U1086 ( .IN1(n1859), .IN2(n1847), .IN3(\mem[25][21] ), .IN4(n1936), 
        .Q(n935) );
  AND2X1 U1087 ( .IN1(wr_data[21]), .IN2(n1837), .Q(n47) );
  AO22X1 U1088 ( .IN1(n1857), .IN2(n1846), .IN3(\mem[25][22] ), .IN4(n1936), 
        .Q(n936) );
  AND2X1 U1089 ( .IN1(wr_data[22]), .IN2(n1836), .Q(n48) );
  AO22X1 U1090 ( .IN1(n1855), .IN2(n113), .IN3(\mem[25][23] ), .IN4(n1936), 
        .Q(n937) );
  AND2X1 U1091 ( .IN1(wr_data[23]), .IN2(n1835), .Q(n49) );
  AO22X1 U1092 ( .IN1(n1854), .IN2(n1847), .IN3(\mem[25][24] ), .IN4(n1936), 
        .Q(n938) );
  AO22X1 U1094 ( .IN1(n1853), .IN2(n1846), .IN3(\mem[25][25] ), .IN4(n1936), 
        .Q(n939) );
  AO22X1 U1096 ( .IN1(n1852), .IN2(n1847), .IN3(\mem[25][26] ), .IN4(n1935), 
        .Q(n940) );
  AO22X1 U1098 ( .IN1(n1851), .IN2(n1846), .IN3(\mem[25][27] ), .IN4(n1936), 
        .Q(n941) );
  AO22X1 U1100 ( .IN1(n1850), .IN2(n1847), .IN3(\mem[25][28] ), .IN4(n1935), 
        .Q(n942) );
  AO22X1 U1102 ( .IN1(n1849), .IN2(n1846), .IN3(\mem[25][29] ), .IN4(n1936), 
        .Q(n943) );
  AO22X1 U1104 ( .IN1(n1848), .IN2(n1847), .IN3(\mem[25][30] ), .IN4(n1935), 
        .Q(n944) );
  AO22X1 U1106 ( .IN1(n1845), .IN2(n1846), .IN3(\mem[25][31] ), .IN4(n1935), 
        .Q(n945) );
  AO21X1 U1107 ( .IN1(n83), .IN2(n73), .IN3(n1999), .Q(n113) );
  AND3X1 U1108 ( .IN1(n2003), .IN2(n2002), .IN3(wr_addr[0]), .Q(n83) );
  AO22X1 U1110 ( .IN1(n1844), .IN2(n1841), .IN3(\mem[26][0] ), .IN4(n1996), 
        .Q(n946) );
  AO22X1 U1112 ( .IN1(n1843), .IN2(n39), .IN3(\mem[26][1] ), .IN4(n1996), .Q(
        n947) );
  AO22X1 U1114 ( .IN1(n61), .IN2(n1842), .IN3(\mem[26][2] ), .IN4(n1996), .Q(
        n948) );
  AO22X1 U1116 ( .IN1(n62), .IN2(n1841), .IN3(\mem[26][3] ), .IN4(n1996), .Q(
        n949) );
  AO22X1 U1118 ( .IN1(n63), .IN2(n39), .IN3(\mem[26][4] ), .IN4(n1996), .Q(
        n950) );
  AO22X1 U1120 ( .IN1(n64), .IN2(n1842), .IN3(\mem[26][5] ), .IN4(n1995), .Q(
        n951) );
  AO22X1 U1122 ( .IN1(n65), .IN2(n1841), .IN3(\mem[26][6] ), .IN4(n1996), .Q(
        n952) );
  AO22X1 U1124 ( .IN1(n66), .IN2(n1842), .IN3(\mem[26][7] ), .IN4(n1996), .Q(
        n953) );
  AO22X1 U1126 ( .IN1(n67), .IN2(n1841), .IN3(\mem[26][8] ), .IN4(n1995), .Q(
        n954) );
  AO22X1 U1128 ( .IN1(n68), .IN2(n1842), .IN3(\mem[26][9] ), .IN4(n1996), .Q(
        n955) );
  AO22X1 U1130 ( .IN1(n69), .IN2(n1841), .IN3(\mem[26][10] ), .IN4(n1995), .Q(
        n956) );
  AO22X1 U1132 ( .IN1(n70), .IN2(n1842), .IN3(\mem[26][11] ), .IN4(n1996), .Q(
        n957) );
  AO22X1 U1134 ( .IN1(n71), .IN2(n1841), .IN3(\mem[26][12] ), .IN4(n1995), .Q(
        n958) );
  AO21X1 U1135 ( .IN1(n86), .IN2(n73), .IN3(n1999), .Q(n39) );
  AND3X1 U1136 ( .IN1(wr_addr[3]), .IN2(n1834), .IN3(wr_addr[4]), .Q(n73) );
  AND3X1 U1137 ( .IN1(n2004), .IN2(n2002), .IN3(wr_addr[1]), .Q(n86) );
  NAND2X1 U3 ( .IN1(wr_en), .IN2(nrst), .QN(n1) );
  AO21X1 U4 ( .IN1(n104), .IN2(n72), .IN3(n1998), .Q(n107) );
  AO21X1 U5 ( .IN1(n104), .IN2(n86), .IN3(n1998), .Q(n106) );
  AO21X1 U6 ( .IN1(n104), .IN2(n83), .IN3(n1998), .Q(n105) );
  AO21X1 U7 ( .IN1(n104), .IN2(n94), .IN3(n1998), .Q(n103) );
  AO21X1 U8 ( .IN1(n95), .IN2(n72), .IN3(n1998), .Q(n98) );
  AO21X1 U9 ( .IN1(n95), .IN2(n86), .IN3(n1998), .Q(n97) );
  AO21X1 U10 ( .IN1(n95), .IN2(n83), .IN3(n1998), .Q(n96) );
  AO21X1 U11 ( .IN1(n94), .IN2(n95), .IN3(n1998), .Q(n93) );
  AO21X1 U12 ( .IN1(n84), .IN2(n77), .IN3(n1997), .Q(n89) );
  AO21X1 U13 ( .IN1(n84), .IN2(n75), .IN3(n1997), .Q(n88) );
  AO21X1 U14 ( .IN1(n84), .IN2(n72), .IN3(n1997), .Q(n87) );
  AO21X1 U15 ( .IN1(n84), .IN2(n86), .IN3(n1997), .Q(n85) );
  AO21X1 U16 ( .IN1(n83), .IN2(n84), .IN3(n1997), .Q(n82) );
  AO21X1 U17 ( .IN1(n81), .IN2(n73), .IN3(n1997), .Q(n80) );
  AO21X1 U18 ( .IN1(n79), .IN2(n73), .IN3(n1997), .Q(n78) );
  AO21X1 U19 ( .IN1(n77), .IN2(n73), .IN3(n1997), .Q(n76) );
  AO21X1 U20 ( .IN1(n75), .IN2(n73), .IN3(n1997), .Q(n74) );
  AO21X1 U21 ( .IN1(n72), .IN2(n73), .IN3(n1997), .Q(n59) );
  INVX0 U22 ( .INP(N11), .ZN(n1427) );
  INVX0 U23 ( .INP(N10), .ZN(n1446) );
  INVX0 U24 ( .INP(N15), .ZN(n1813) );
  INVX0 U25 ( .INP(N16), .ZN(n1792) );
  INVX0 U26 ( .INP(N11), .ZN(n1426) );
  INVX0 U27 ( .INP(N10), .ZN(n1445) );
  INVX0 U28 ( .INP(N15), .ZN(n1812) );
  INVX0 U29 ( .INP(N16), .ZN(n1791) );
  INVX0 U30 ( .INP(N17), .ZN(n1786) );
  INVX0 U31 ( .INP(N12), .ZN(n1421) );
  INVX0 U32 ( .INP(n103), .ZN(n1953) );
  INVX0 U33 ( .INP(n103), .ZN(n1954) );
  INVX0 U34 ( .INP(n105), .ZN(n1951) );
  INVX0 U35 ( .INP(n105), .ZN(n1952) );
  INVX0 U36 ( .INP(n106), .ZN(n1949) );
  INVX0 U37 ( .INP(n106), .ZN(n1950) );
  INVX0 U38 ( .INP(n107), .ZN(n1947) );
  INVX0 U39 ( .INP(n107), .ZN(n1948) );
  INVX0 U91 ( .INP(n96), .ZN(n1967) );
  INVX0 U124 ( .INP(n96), .ZN(n1968) );
  INVX0 U157 ( .INP(n97), .ZN(n1965) );
  INVX0 U190 ( .INP(n97), .ZN(n1966) );
  INVX0 U223 ( .INP(n98), .ZN(n1963) );
  INVX0 U288 ( .INP(n98), .ZN(n1964) );
  INVX0 U321 ( .INP(n85), .ZN(n1981) );
  INVX0 U354 ( .INP(n85), .ZN(n1982) );
  INVX0 U387 ( .INP(n87), .ZN(n1979) );
  INVX0 U420 ( .INP(n87), .ZN(n1980) );
  INVX0 U520 ( .INP(n88), .ZN(n1977) );
  INVX0 U553 ( .INP(n88), .ZN(n1978) );
  INVX0 U586 ( .INP(n89), .ZN(n1975) );
  INVX0 U619 ( .INP(n89), .ZN(n1976) );
  INVX0 U785 ( .INP(n82), .ZN(n1983) );
  INVX0 U818 ( .INP(n82), .ZN(n1984) );
  INVX0 U851 ( .INP(n59), .ZN(n1993) );
  INVX0 U884 ( .INP(n59), .ZN(n1994) );
  INVX0 U1071 ( .INP(n74), .ZN(n1991) );
  INVX0 U1073 ( .INP(n74), .ZN(n1992) );
  INVX0 U1075 ( .INP(n76), .ZN(n1989) );
  INVX0 U1093 ( .INP(n76), .ZN(n1990) );
  INVX0 U1095 ( .INP(n78), .ZN(n1987) );
  INVX0 U1097 ( .INP(n78), .ZN(n1988) );
  INVX0 U1099 ( .INP(n80), .ZN(n1985) );
  INVX0 U1101 ( .INP(n80), .ZN(n1986) );
  INVX0 U1103 ( .INP(n93), .ZN(n1969) );
  INVX0 U1105 ( .INP(n93), .ZN(n1970) );
  INVX0 U1109 ( .INP(n112), .ZN(n1937) );
  INVX0 U1111 ( .INP(n112), .ZN(n1938) );
  INVX0 U1113 ( .INP(n113), .ZN(n1935) );
  INVX0 U1115 ( .INP(n113), .ZN(n1936) );
  INVX0 U1117 ( .INP(n39), .ZN(n1995) );
  INVX0 U1119 ( .INP(n39), .ZN(n1996) );
  INVX0 U1121 ( .INP(n90), .ZN(n1973) );
  INVX0 U1123 ( .INP(n90), .ZN(n1974) );
  INVX0 U1125 ( .INP(n91), .ZN(n1971) );
  INVX0 U1127 ( .INP(n91), .ZN(n1972) );
  INVX0 U1129 ( .INP(n99), .ZN(n1961) );
  INVX0 U1131 ( .INP(n99), .ZN(n1962) );
  INVX0 U1133 ( .INP(n100), .ZN(n1959) );
  INVX0 U1138 ( .INP(n100), .ZN(n1960) );
  INVX0 U1139 ( .INP(n101), .ZN(n1957) );
  INVX0 U1140 ( .INP(n101), .ZN(n1958) );
  INVX0 U1141 ( .INP(n102), .ZN(n1955) );
  INVX0 U1142 ( .INP(n102), .ZN(n1956) );
  INVX0 U1143 ( .INP(n108), .ZN(n1945) );
  INVX0 U1144 ( .INP(n108), .ZN(n1946) );
  INVX0 U1145 ( .INP(n109), .ZN(n1943) );
  INVX0 U1146 ( .INP(n109), .ZN(n1944) );
  INVX0 U1147 ( .INP(n110), .ZN(n1941) );
  INVX0 U1148 ( .INP(n110), .ZN(n1942) );
  INVX0 U1149 ( .INP(n111), .ZN(n1939) );
  INVX0 U1150 ( .INP(n111), .ZN(n1940) );
  INVX0 U1151 ( .INP(n1), .ZN(n1838) );
  INVX0 U1152 ( .INP(n1), .ZN(n1834) );
  INVX0 U1153 ( .INP(n1), .ZN(n1836) );
  INVX0 U1154 ( .INP(n1), .ZN(n1835) );
  INVX0 U1155 ( .INP(n1), .ZN(n1837) );
  INVX0 U1156 ( .INP(n1), .ZN(n1840) );
  INVX0 U1157 ( .INP(n1), .ZN(n1839) );
  INVX0 U1158 ( .INP(n1813), .ZN(n1814) );
  INVX0 U1159 ( .INP(n1813), .ZN(n1815) );
  INVX0 U1160 ( .INP(n1813), .ZN(n1816) );
  INVX0 U1161 ( .INP(n1813), .ZN(n1817) );
  INVX0 U1162 ( .INP(n1813), .ZN(n1818) );
  INVX0 U1163 ( .INP(n1813), .ZN(n1819) );
  INVX0 U1164 ( .INP(n1813), .ZN(n1820) );
  INVX0 U1165 ( .INP(n1813), .ZN(n1821) );
  INVX0 U1166 ( .INP(n1813), .ZN(n1822) );
  INVX0 U1167 ( .INP(n1813), .ZN(n1823) );
  INVX0 U1168 ( .INP(n1813), .ZN(n1824) );
  INVX0 U1169 ( .INP(n1446), .ZN(n1447) );
  INVX0 U1170 ( .INP(n1446), .ZN(n1448) );
  INVX0 U1171 ( .INP(n1446), .ZN(n1449) );
  INVX0 U1172 ( .INP(n1446), .ZN(n1450) );
  INVX0 U1173 ( .INP(n1446), .ZN(n1451) );
  INVX0 U1174 ( .INP(n1446), .ZN(n1452) );
  INVX0 U1175 ( .INP(n1446), .ZN(n1453) );
  INVX0 U1176 ( .INP(n1446), .ZN(n1454) );
  INVX0 U1177 ( .INP(n1446), .ZN(n1455) );
  INVX0 U1178 ( .INP(n1446), .ZN(n1456) );
  INVX0 U1179 ( .INP(n1792), .ZN(n1793) );
  INVX0 U1180 ( .INP(n1792), .ZN(n1794) );
  INVX0 U1181 ( .INP(n1792), .ZN(n1795) );
  INVX0 U1182 ( .INP(n1792), .ZN(n1796) );
  INVX0 U1183 ( .INP(n1792), .ZN(n1797) );
  INVX0 U1184 ( .INP(n1792), .ZN(n1798) );
  INVX0 U1185 ( .INP(n1792), .ZN(n1799) );
  INVX0 U1186 ( .INP(n1792), .ZN(n1800) );
  INVX0 U1187 ( .INP(n1792), .ZN(n1801) );
  INVX0 U1188 ( .INP(n1792), .ZN(n1802) );
  INVX0 U1189 ( .INP(n1427), .ZN(n1428) );
  INVX0 U1190 ( .INP(n1427), .ZN(n1429) );
  INVX0 U1191 ( .INP(n1427), .ZN(n1430) );
  INVX0 U1192 ( .INP(n1427), .ZN(n1431) );
  INVX0 U1193 ( .INP(n1427), .ZN(n1432) );
  INVX0 U1194 ( .INP(n1427), .ZN(n1433) );
  INVX0 U1195 ( .INP(n1427), .ZN(n1434) );
  INVX0 U1196 ( .INP(n1427), .ZN(n1435) );
  INVX0 U1197 ( .INP(n1427), .ZN(n1436) );
  INVX0 U1198 ( .INP(n1812), .ZN(n1825) );
  INVX0 U1199 ( .INP(n1812), .ZN(n1826) );
  INVX0 U1200 ( .INP(n1812), .ZN(n1827) );
  INVX0 U1201 ( .INP(n1812), .ZN(n1828) );
  INVX0 U1202 ( .INP(n1812), .ZN(n1829) );
  INVX0 U1203 ( .INP(n1812), .ZN(n1830) );
  INVX0 U1204 ( .INP(n1812), .ZN(n1831) );
  INVX0 U1205 ( .INP(n1812), .ZN(n1832) );
  INVX0 U1206 ( .INP(n1812), .ZN(n1833) );
  INVX0 U1207 ( .INP(n1445), .ZN(n1457) );
  INVX0 U1208 ( .INP(n1445), .ZN(n1458) );
  INVX0 U1209 ( .INP(n1445), .ZN(n1459) );
  INVX0 U1210 ( .INP(n1445), .ZN(n1460) );
  INVX0 U1211 ( .INP(n1445), .ZN(n1461) );
  INVX0 U1212 ( .INP(n1445), .ZN(n1462) );
  INVX0 U1213 ( .INP(n1445), .ZN(n1463) );
  INVX0 U1214 ( .INP(n1445), .ZN(n1464) );
  INVX0 U1215 ( .INP(n1445), .ZN(n1465) );
  INVX0 U1216 ( .INP(n1791), .ZN(n1803) );
  INVX0 U1217 ( .INP(n1791), .ZN(n1804) );
  INVX0 U1218 ( .INP(n1791), .ZN(n1805) );
  INVX0 U1219 ( .INP(n1791), .ZN(n1806) );
  INVX0 U1220 ( .INP(n1791), .ZN(n1807) );
  INVX0 U1221 ( .INP(n1791), .ZN(n1808) );
  INVX0 U1222 ( .INP(n1791), .ZN(n1809) );
  INVX0 U1223 ( .INP(n1791), .ZN(n1810) );
  INVX0 U1224 ( .INP(n1791), .ZN(n1811) );
  INVX0 U1225 ( .INP(n1426), .ZN(n1437) );
  INVX0 U1226 ( .INP(n1426), .ZN(n1438) );
  INVX0 U1227 ( .INP(n1426), .ZN(n1439) );
  INVX0 U1228 ( .INP(n1426), .ZN(n1440) );
  INVX0 U1229 ( .INP(n1426), .ZN(n1441) );
  INVX0 U1230 ( .INP(n1426), .ZN(n1442) );
  INVX0 U1231 ( .INP(n1426), .ZN(n1443) );
  INVX0 U1232 ( .INP(n1426), .ZN(n1444) );
  INVX0 U1233 ( .INP(n1786), .ZN(n1790) );
  INVX0 U1234 ( .INP(n1786), .ZN(n1789) );
  INVX0 U1235 ( .INP(n1786), .ZN(n1788) );
  INVX0 U1236 ( .INP(n1421), .ZN(n1425) );
  INVX0 U1237 ( .INP(n1421), .ZN(n1424) );
  INVX0 U1238 ( .INP(n1786), .ZN(n1787) );
  INVX0 U1239 ( .INP(n1421), .ZN(n1423) );
  INVX0 U1240 ( .INP(n1421), .ZN(n1422) );
  AO21X1 U1241 ( .IN1(n104), .IN2(n94), .IN3(n1998), .Q(n1894) );
  AO21X1 U1242 ( .IN1(n104), .IN2(n94), .IN3(n1998), .Q(n1893) );
  AO21X1 U1243 ( .IN1(n104), .IN2(n83), .IN3(n1998), .Q(n1892) );
  AO21X1 U1244 ( .IN1(n104), .IN2(n83), .IN3(n1998), .Q(n1891) );
  AO21X1 U1245 ( .IN1(n104), .IN2(n86), .IN3(n1998), .Q(n1890) );
  AO21X1 U1246 ( .IN1(n104), .IN2(n86), .IN3(n1998), .Q(n1889) );
  AO21X1 U1247 ( .IN1(n104), .IN2(n72), .IN3(n1998), .Q(n1888) );
  AO21X1 U1248 ( .IN1(n104), .IN2(n72), .IN3(n1998), .Q(n1887) );
  AO21X1 U1249 ( .IN1(n95), .IN2(n83), .IN3(n1998), .Q(n1908) );
  AO21X1 U1250 ( .IN1(n95), .IN2(n83), .IN3(n1998), .Q(n1907) );
  AO21X1 U1251 ( .IN1(n95), .IN2(n86), .IN3(n1998), .Q(n1906) );
  AO21X1 U1252 ( .IN1(n95), .IN2(n86), .IN3(n1998), .Q(n1905) );
  AO21X1 U1253 ( .IN1(n95), .IN2(n72), .IN3(n1998), .Q(n1904) );
  AO21X1 U1254 ( .IN1(n95), .IN2(n72), .IN3(n1998), .Q(n1903) );
  AO21X1 U1255 ( .IN1(n84), .IN2(n86), .IN3(n1997), .Q(n1922) );
  AO21X1 U1256 ( .IN1(n84), .IN2(n86), .IN3(n1997), .Q(n1921) );
  AO21X1 U1257 ( .IN1(n84), .IN2(n72), .IN3(n1997), .Q(n1920) );
  AO21X1 U1258 ( .IN1(n84), .IN2(n72), .IN3(n1997), .Q(n1919) );
  AO21X1 U1259 ( .IN1(n84), .IN2(n75), .IN3(n1997), .Q(n1918) );
  AO21X1 U1260 ( .IN1(n84), .IN2(n75), .IN3(n1997), .Q(n1917) );
  AO21X1 U1261 ( .IN1(n94), .IN2(n95), .IN3(n1998), .Q(n1910) );
  AO21X1 U1262 ( .IN1(n94), .IN2(n95), .IN3(n1998), .Q(n1909) );
  AO21X1 U1263 ( .IN1(n72), .IN2(n73), .IN3(n1997), .Q(n1934) );
  AO21X1 U1264 ( .IN1(n72), .IN2(n73), .IN3(n1997), .Q(n1933) );
  AO21X1 U1265 ( .IN1(n75), .IN2(n73), .IN3(n1997), .Q(n1932) );
  AO21X1 U1266 ( .IN1(n75), .IN2(n73), .IN3(n1997), .Q(n1931) );
  AO21X1 U1267 ( .IN1(n77), .IN2(n73), .IN3(n1997), .Q(n1930) );
  AO21X1 U1268 ( .IN1(n77), .IN2(n73), .IN3(n1997), .Q(n1929) );
  AO21X1 U1269 ( .IN1(n79), .IN2(n73), .IN3(n1997), .Q(n1928) );
  AO21X1 U1270 ( .IN1(n79), .IN2(n73), .IN3(n1997), .Q(n1927) );
  AO21X1 U1271 ( .IN1(n83), .IN2(n84), .IN3(n1997), .Q(n1924) );
  AO21X1 U1272 ( .IN1(n83), .IN2(n84), .IN3(n1997), .Q(n1923) );
  AND2X1 U1273 ( .IN1(wr_data[3]), .IN2(n1838), .Q(n62) );
  AND2X1 U1274 ( .IN1(wr_data[5]), .IN2(n1838), .Q(n64) );
  AND2X1 U1275 ( .IN1(wr_data[10]), .IN2(n1838), .Q(n69) );
  AND2X1 U1276 ( .IN1(wr_data[2]), .IN2(n1835), .Q(n61) );
  AND2X1 U1277 ( .IN1(wr_data[4]), .IN2(n1836), .Q(n63) );
  AND2X1 U1278 ( .IN1(wr_data[11]), .IN2(n1834), .Q(n70) );
  AND2X1 U1279 ( .IN1(wr_data[6]), .IN2(n1837), .Q(n65) );
  AND2X1 U1280 ( .IN1(wr_data[12]), .IN2(n1837), .Q(n71) );
  AND2X1 U1281 ( .IN1(wr_data[7]), .IN2(n1839), .Q(n66) );
  AND2X1 U1282 ( .IN1(wr_data[8]), .IN2(n1839), .Q(n67) );
  AND2X1 U1283 ( .IN1(wr_data[9]), .IN2(n1839), .Q(n68) );
  INVX0 U1284 ( .INP(nrst), .ZN(n1998) );
  INVX0 U1285 ( .INP(nrst), .ZN(n1997) );
  INVX0 U1286 ( .INP(nrst), .ZN(n1999) );
  AND2X1 U1287 ( .IN1(wr_data[25]), .IN2(n1840), .Q(n1853) );
  AND2X1 U1288 ( .IN1(wr_data[26]), .IN2(n1840), .Q(n1852) );
  AND2X1 U1289 ( .IN1(wr_data[27]), .IN2(n1840), .Q(n1851) );
  AND2X1 U1290 ( .IN1(wr_data[28]), .IN2(n1836), .Q(n1850) );
  AND2X1 U1291 ( .IN1(wr_data[29]), .IN2(n1836), .Q(n1849) );
  AND2X1 U1292 ( .IN1(wr_data[30]), .IN2(n1837), .Q(n1848) );
  AND2X1 U1293 ( .IN1(wr_data[31]), .IN2(n1839), .Q(n1845) );
  AND2X1 U1294 ( .IN1(wr_data[24]), .IN2(n1838), .Q(n1854) );
  AND2X1 U1295 ( .IN1(wr_data[0]), .IN2(n1834), .Q(n1844) );
  AND2X1 U1296 ( .IN1(wr_data[1]), .IN2(n1840), .Q(n1843) );
  AND2X1 U1297 ( .IN1(wr_data[25]), .IN2(n1837), .Q(n51) );
  AND2X1 U1298 ( .IN1(wr_data[26]), .IN2(n1838), .Q(n52) );
  AND2X1 U1299 ( .IN1(wr_data[27]), .IN2(n1840), .Q(n53) );
  AND2X1 U1300 ( .IN1(wr_data[28]), .IN2(n1837), .Q(n54) );
  AND2X1 U1301 ( .IN1(wr_data[29]), .IN2(n1835), .Q(n55) );
  AND2X1 U1302 ( .IN1(wr_data[30]), .IN2(n1839), .Q(n56) );
  AND2X1 U1303 ( .IN1(wr_data[31]), .IN2(n1840), .Q(n57) );
  AND2X1 U1304 ( .IN1(wr_data[0]), .IN2(n1840), .Q(n58) );
  AND2X1 U1305 ( .IN1(wr_data[1]), .IN2(n1840), .Q(n60) );
  AND2X1 U1306 ( .IN1(wr_data[24]), .IN2(n1839), .Q(n50) );
  AND2X1 U1307 ( .IN1(wr_data[13]), .IN2(n1840), .Q(n1875) );
  AND2X1 U1308 ( .IN1(wr_data[14]), .IN2(n1835), .Q(n40) );
  AND2X1 U1309 ( .IN1(wr_data[15]), .IN2(n1840), .Q(n41) );
  AND2X1 U1310 ( .IN1(wr_data[14]), .IN2(n1834), .Q(n1874) );
  AND2X1 U1311 ( .IN1(wr_data[15]), .IN2(n1839), .Q(n1872) );
  AND2X1 U1312 ( .IN1(wr_data[13]), .IN2(n1838), .Q(n38) );
  AND2X1 U1313 ( .IN1(wr_data[13]), .IN2(n1839), .Q(n1876) );
  INVX0 U1314 ( .INP(wr_addr[2]), .ZN(n2002) );
  INVX0 U1315 ( .INP(wr_addr[1]), .ZN(n2003) );
  INVX0 U1316 ( .INP(wr_addr[0]), .ZN(n2004) );
  INVX0 U1317 ( .INP(wr_addr[4]), .ZN(n2000) );
  INVX0 U1318 ( .INP(wr_addr[3]), .ZN(n2001) );
  MUX41X1 U1319 ( .IN1(\mem[28][0] ), .IN3(\mem[30][0] ), .IN2(\mem[29][0] ), 
        .IN4(\mem[31][0] ), .S0(n1439), .S1(N10), .Q(n2) );
  MUX41X1 U1320 ( .IN1(\mem[24][0] ), .IN3(\mem[26][0] ), .IN2(\mem[25][0] ), 
        .IN4(\mem[27][0] ), .S0(n1438), .S1(N10), .Q(n3) );
  MUX41X1 U1321 ( .IN1(\mem[20][0] ), .IN3(\mem[22][0] ), .IN2(\mem[21][0] ), 
        .IN4(\mem[23][0] ), .S0(n1437), .S1(N10), .Q(n4) );
  MUX41X1 U1322 ( .IN1(\mem[16][0] ), .IN3(\mem[18][0] ), .IN2(\mem[17][0] ), 
        .IN4(\mem[19][0] ), .S0(n1438), .S1(n1463), .Q(n5) );
  MUX41X1 U1323 ( .IN1(n5), .IN3(n3), .IN2(n4), .IN4(n2), .S0(N13), .S1(n1425), 
        .Q(n6) );
  MUX41X1 U1324 ( .IN1(\mem[12][0] ), .IN3(\mem[14][0] ), .IN2(\mem[13][0] ), 
        .IN4(\mem[15][0] ), .S0(n1428), .S1(n1447), .Q(n7) );
  MUX41X1 U1325 ( .IN1(\mem[8][0] ), .IN3(\mem[10][0] ), .IN2(\mem[9][0] ), 
        .IN4(\mem[11][0] ), .S0(n1428), .S1(n1447), .Q(n8) );
  MUX41X1 U1326 ( .IN1(\mem[4][0] ), .IN3(\mem[6][0] ), .IN2(\mem[5][0] ), 
        .IN4(\mem[7][0] ), .S0(n1428), .S1(n1447), .Q(n9) );
  MUX41X1 U1327 ( .IN1(\mem[0][0] ), .IN3(\mem[2][0] ), .IN2(\mem[1][0] ), 
        .IN4(\mem[3][0] ), .S0(n1428), .S1(n1447), .Q(n10) );
  MUX41X1 U1328 ( .IN1(n10), .IN3(n8), .IN2(n9), .IN4(n7), .S0(N13), .S1(n1425), .Q(n11) );
  MUX21X1 U1329 ( .IN1(n11), .IN2(n6), .S(N14), .Q(rd_dataA[0]) );
  MUX41X1 U1330 ( .IN1(\mem[28][1] ), .IN3(\mem[30][1] ), .IN2(\mem[29][1] ), 
        .IN4(\mem[31][1] ), .S0(n1428), .S1(n1447), .Q(n12) );
  MUX41X1 U1331 ( .IN1(\mem[24][1] ), .IN3(\mem[26][1] ), .IN2(\mem[25][1] ), 
        .IN4(\mem[27][1] ), .S0(n1428), .S1(n1447), .Q(n13) );
  MUX41X1 U1332 ( .IN1(\mem[20][1] ), .IN3(\mem[22][1] ), .IN2(\mem[21][1] ), 
        .IN4(\mem[23][1] ), .S0(n1428), .S1(n1447), .Q(n14) );
  MUX41X1 U1333 ( .IN1(\mem[16][1] ), .IN3(\mem[18][1] ), .IN2(\mem[17][1] ), 
        .IN4(\mem[19][1] ), .S0(n1428), .S1(n1447), .Q(n15) );
  MUX41X1 U1334 ( .IN1(n15), .IN3(n13), .IN2(n14), .IN4(n12), .S0(N13), .S1(
        n1425), .Q(n16) );
  MUX41X1 U1335 ( .IN1(\mem[12][1] ), .IN3(\mem[14][1] ), .IN2(\mem[13][1] ), 
        .IN4(\mem[15][1] ), .S0(n1428), .S1(n1447), .Q(n17) );
  MUX41X1 U1336 ( .IN1(\mem[8][1] ), .IN3(\mem[10][1] ), .IN2(\mem[9][1] ), 
        .IN4(\mem[11][1] ), .S0(n1428), .S1(n1447), .Q(n18) );
  MUX41X1 U1337 ( .IN1(\mem[4][1] ), .IN3(\mem[6][1] ), .IN2(\mem[5][1] ), 
        .IN4(\mem[7][1] ), .S0(n1428), .S1(n1447), .Q(n19) );
  MUX41X1 U1338 ( .IN1(\mem[0][1] ), .IN3(\mem[2][1] ), .IN2(\mem[1][1] ), 
        .IN4(\mem[3][1] ), .S0(n1428), .S1(n1447), .Q(n20) );
  MUX41X1 U1339 ( .IN1(n20), .IN3(n18), .IN2(n19), .IN4(n17), .S0(N13), .S1(
        n1425), .Q(n21) );
  MUX21X1 U1340 ( .IN1(n21), .IN2(n16), .S(N14), .Q(rd_dataA[1]) );
  MUX41X1 U1341 ( .IN1(\mem[28][2] ), .IN3(\mem[30][2] ), .IN2(\mem[29][2] ), 
        .IN4(\mem[31][2] ), .S0(n1429), .S1(n1448), .Q(n22) );
  MUX41X1 U1342 ( .IN1(\mem[24][2] ), .IN3(\mem[26][2] ), .IN2(\mem[25][2] ), 
        .IN4(\mem[27][2] ), .S0(n1429), .S1(n1448), .Q(n23) );
  MUX41X1 U1343 ( .IN1(\mem[20][2] ), .IN3(\mem[22][2] ), .IN2(\mem[21][2] ), 
        .IN4(\mem[23][2] ), .S0(n1429), .S1(n1448), .Q(n24) );
  MUX41X1 U1344 ( .IN1(\mem[16][2] ), .IN3(\mem[18][2] ), .IN2(\mem[17][2] ), 
        .IN4(\mem[19][2] ), .S0(n1429), .S1(n1448), .Q(n25) );
  MUX41X1 U1345 ( .IN1(n25), .IN3(n23), .IN2(n24), .IN4(n22), .S0(N13), .S1(
        n1425), .Q(n26) );
  MUX41X1 U1346 ( .IN1(\mem[12][2] ), .IN3(\mem[14][2] ), .IN2(\mem[13][2] ), 
        .IN4(\mem[15][2] ), .S0(n1429), .S1(n1448), .Q(n27) );
  MUX41X1 U1347 ( .IN1(\mem[8][2] ), .IN3(\mem[10][2] ), .IN2(\mem[9][2] ), 
        .IN4(\mem[11][2] ), .S0(n1429), .S1(n1448), .Q(n28) );
  MUX41X1 U1348 ( .IN1(\mem[4][2] ), .IN3(\mem[6][2] ), .IN2(\mem[5][2] ), 
        .IN4(\mem[7][2] ), .S0(n1429), .S1(n1448), .Q(n29) );
  MUX41X1 U1349 ( .IN1(\mem[0][2] ), .IN3(\mem[2][2] ), .IN2(\mem[1][2] ), 
        .IN4(\mem[3][2] ), .S0(n1429), .S1(n1448), .Q(n30) );
  MUX41X1 U1350 ( .IN1(n30), .IN3(n28), .IN2(n29), .IN4(n27), .S0(N13), .S1(
        n1425), .Q(n31) );
  MUX21X1 U1351 ( .IN1(n31), .IN2(n26), .S(N14), .Q(rd_dataA[2]) );
  MUX41X1 U1352 ( .IN1(\mem[28][3] ), .IN3(\mem[30][3] ), .IN2(\mem[29][3] ), 
        .IN4(\mem[31][3] ), .S0(n1429), .S1(n1448), .Q(n32) );
  MUX41X1 U1353 ( .IN1(\mem[24][3] ), .IN3(\mem[26][3] ), .IN2(\mem[25][3] ), 
        .IN4(\mem[27][3] ), .S0(n1429), .S1(n1448), .Q(n33) );
  MUX41X1 U1354 ( .IN1(\mem[20][3] ), .IN3(\mem[22][3] ), .IN2(\mem[21][3] ), 
        .IN4(\mem[23][3] ), .S0(n1429), .S1(n1448), .Q(n34) );
  MUX41X1 U1355 ( .IN1(\mem[16][3] ), .IN3(\mem[18][3] ), .IN2(\mem[17][3] ), 
        .IN4(\mem[19][3] ), .S0(n1429), .S1(n1448), .Q(n35) );
  MUX41X1 U1356 ( .IN1(n35), .IN3(n33), .IN2(n34), .IN4(n32), .S0(N13), .S1(
        n1425), .Q(n36) );
  MUX41X1 U1357 ( .IN1(\mem[12][3] ), .IN3(\mem[14][3] ), .IN2(\mem[13][3] ), 
        .IN4(\mem[15][3] ), .S0(n1430), .S1(n1449), .Q(n37) );
  MUX41X1 U1358 ( .IN1(\mem[8][3] ), .IN3(\mem[10][3] ), .IN2(\mem[9][3] ), 
        .IN4(\mem[11][3] ), .S0(n1430), .S1(n1449), .Q(n92) );
  MUX41X1 U1359 ( .IN1(\mem[4][3] ), .IN3(\mem[6][3] ), .IN2(\mem[5][3] ), 
        .IN4(\mem[7][3] ), .S0(n1430), .S1(n1449), .Q(n1138) );
  MUX41X1 U1360 ( .IN1(\mem[0][3] ), .IN3(\mem[2][3] ), .IN2(\mem[1][3] ), 
        .IN4(\mem[3][3] ), .S0(n1430), .S1(n1449), .Q(n1139) );
  MUX41X1 U1361 ( .IN1(n1139), .IN3(n92), .IN2(n1138), .IN4(n37), .S0(N13), 
        .S1(n1425), .Q(n1140) );
  MUX21X1 U1362 ( .IN1(n1140), .IN2(n36), .S(N14), .Q(rd_dataA[3]) );
  MUX41X1 U1363 ( .IN1(\mem[28][4] ), .IN3(\mem[30][4] ), .IN2(\mem[29][4] ), 
        .IN4(\mem[31][4] ), .S0(n1430), .S1(n1449), .Q(n1141) );
  MUX41X1 U1364 ( .IN1(\mem[24][4] ), .IN3(\mem[26][4] ), .IN2(\mem[25][4] ), 
        .IN4(\mem[27][4] ), .S0(n1430), .S1(n1449), .Q(n1142) );
  MUX41X1 U1365 ( .IN1(\mem[20][4] ), .IN3(\mem[22][4] ), .IN2(\mem[21][4] ), 
        .IN4(\mem[23][4] ), .S0(n1430), .S1(n1449), .Q(n1143) );
  MUX41X1 U1366 ( .IN1(\mem[16][4] ), .IN3(\mem[18][4] ), .IN2(\mem[17][4] ), 
        .IN4(\mem[19][4] ), .S0(n1430), .S1(n1449), .Q(n1144) );
  MUX41X1 U1367 ( .IN1(n1144), .IN3(n1142), .IN2(n1143), .IN4(n1141), .S0(N13), 
        .S1(n1425), .Q(n1145) );
  MUX41X1 U1368 ( .IN1(\mem[12][4] ), .IN3(\mem[14][4] ), .IN2(\mem[13][4] ), 
        .IN4(\mem[15][4] ), .S0(n1430), .S1(n1449), .Q(n1146) );
  MUX41X1 U1369 ( .IN1(\mem[8][4] ), .IN3(\mem[10][4] ), .IN2(\mem[9][4] ), 
        .IN4(\mem[11][4] ), .S0(n1430), .S1(n1449), .Q(n1147) );
  MUX41X1 U1370 ( .IN1(\mem[4][4] ), .IN3(\mem[6][4] ), .IN2(\mem[5][4] ), 
        .IN4(\mem[7][4] ), .S0(n1430), .S1(n1449), .Q(n1148) );
  MUX41X1 U1371 ( .IN1(\mem[0][4] ), .IN3(\mem[2][4] ), .IN2(\mem[1][4] ), 
        .IN4(\mem[3][4] ), .S0(n1430), .S1(n1449), .Q(n1149) );
  MUX41X1 U1372 ( .IN1(n1149), .IN3(n1147), .IN2(n1148), .IN4(n1146), .S0(N13), 
        .S1(n1425), .Q(n1150) );
  MUX21X1 U1373 ( .IN1(n1150), .IN2(n1145), .S(N14), .Q(rd_dataA[4]) );
  MUX41X1 U1374 ( .IN1(\mem[28][5] ), .IN3(\mem[30][5] ), .IN2(\mem[29][5] ), 
        .IN4(\mem[31][5] ), .S0(n1431), .S1(n1450), .Q(n1151) );
  MUX41X1 U1375 ( .IN1(\mem[24][5] ), .IN3(\mem[26][5] ), .IN2(\mem[25][5] ), 
        .IN4(\mem[27][5] ), .S0(n1431), .S1(n1450), .Q(n1152) );
  MUX41X1 U1376 ( .IN1(\mem[20][5] ), .IN3(\mem[22][5] ), .IN2(\mem[21][5] ), 
        .IN4(\mem[23][5] ), .S0(n1431), .S1(n1450), .Q(n1153) );
  MUX41X1 U1377 ( .IN1(\mem[16][5] ), .IN3(\mem[18][5] ), .IN2(\mem[17][5] ), 
        .IN4(\mem[19][5] ), .S0(n1431), .S1(n1450), .Q(n1154) );
  MUX41X1 U1378 ( .IN1(n1154), .IN3(n1152), .IN2(n1153), .IN4(n1151), .S0(N13), 
        .S1(n1425), .Q(n1155) );
  MUX41X1 U1379 ( .IN1(\mem[12][5] ), .IN3(\mem[14][5] ), .IN2(\mem[13][5] ), 
        .IN4(\mem[15][5] ), .S0(n1431), .S1(n1450), .Q(n1156) );
  MUX41X1 U1380 ( .IN1(\mem[8][5] ), .IN3(\mem[10][5] ), .IN2(\mem[9][5] ), 
        .IN4(\mem[11][5] ), .S0(n1431), .S1(n1450), .Q(n1157) );
  MUX41X1 U1381 ( .IN1(\mem[4][5] ), .IN3(\mem[6][5] ), .IN2(\mem[5][5] ), 
        .IN4(\mem[7][5] ), .S0(n1431), .S1(n1450), .Q(n1158) );
  MUX41X1 U1382 ( .IN1(\mem[0][5] ), .IN3(\mem[2][5] ), .IN2(\mem[1][5] ), 
        .IN4(\mem[3][5] ), .S0(n1431), .S1(n1450), .Q(n1159) );
  MUX41X1 U1383 ( .IN1(n1159), .IN3(n1157), .IN2(n1158), .IN4(n1156), .S0(N13), 
        .S1(n1425), .Q(n1160) );
  MUX21X1 U1384 ( .IN1(n1160), .IN2(n1155), .S(N14), .Q(rd_dataA[5]) );
  MUX41X1 U1385 ( .IN1(\mem[28][6] ), .IN3(\mem[30][6] ), .IN2(\mem[29][6] ), 
        .IN4(\mem[31][6] ), .S0(n1431), .S1(n1450), .Q(n1161) );
  MUX41X1 U1386 ( .IN1(\mem[24][6] ), .IN3(\mem[26][6] ), .IN2(\mem[25][6] ), 
        .IN4(\mem[27][6] ), .S0(n1431), .S1(n1450), .Q(n1162) );
  MUX41X1 U1387 ( .IN1(\mem[20][6] ), .IN3(\mem[22][6] ), .IN2(\mem[21][6] ), 
        .IN4(\mem[23][6] ), .S0(n1431), .S1(n1450), .Q(n1163) );
  MUX41X1 U1388 ( .IN1(\mem[16][6] ), .IN3(\mem[18][6] ), .IN2(\mem[17][6] ), 
        .IN4(\mem[19][6] ), .S0(n1431), .S1(n1450), .Q(n1164) );
  MUX41X1 U1389 ( .IN1(n1164), .IN3(n1162), .IN2(n1163), .IN4(n1161), .S0(N13), 
        .S1(n1424), .Q(n1165) );
  MUX41X1 U1390 ( .IN1(\mem[12][6] ), .IN3(\mem[14][6] ), .IN2(\mem[13][6] ), 
        .IN4(\mem[15][6] ), .S0(n1432), .S1(n1451), .Q(n1166) );
  MUX41X1 U1391 ( .IN1(\mem[8][6] ), .IN3(\mem[10][6] ), .IN2(\mem[9][6] ), 
        .IN4(\mem[11][6] ), .S0(n1432), .S1(n1451), .Q(n1167) );
  MUX41X1 U1392 ( .IN1(\mem[4][6] ), .IN3(\mem[6][6] ), .IN2(\mem[5][6] ), 
        .IN4(\mem[7][6] ), .S0(n1432), .S1(n1451), .Q(n1168) );
  MUX41X1 U1393 ( .IN1(\mem[0][6] ), .IN3(\mem[2][6] ), .IN2(\mem[1][6] ), 
        .IN4(\mem[3][6] ), .S0(n1432), .S1(n1451), .Q(n1169) );
  MUX41X1 U1394 ( .IN1(n1169), .IN3(n1167), .IN2(n1168), .IN4(n1166), .S0(N13), 
        .S1(n1424), .Q(n1170) );
  MUX21X1 U1395 ( .IN1(n1170), .IN2(n1165), .S(N14), .Q(rd_dataA[6]) );
  MUX41X1 U1396 ( .IN1(\mem[28][7] ), .IN3(\mem[30][7] ), .IN2(\mem[29][7] ), 
        .IN4(\mem[31][7] ), .S0(n1432), .S1(n1451), .Q(n1171) );
  MUX41X1 U1397 ( .IN1(\mem[24][7] ), .IN3(\mem[26][7] ), .IN2(\mem[25][7] ), 
        .IN4(\mem[27][7] ), .S0(n1432), .S1(n1451), .Q(n1172) );
  MUX41X1 U1398 ( .IN1(\mem[20][7] ), .IN3(\mem[22][7] ), .IN2(\mem[21][7] ), 
        .IN4(\mem[23][7] ), .S0(n1432), .S1(n1451), .Q(n1173) );
  MUX41X1 U1399 ( .IN1(\mem[16][7] ), .IN3(\mem[18][7] ), .IN2(\mem[17][7] ), 
        .IN4(\mem[19][7] ), .S0(n1432), .S1(n1451), .Q(n1174) );
  MUX41X1 U1400 ( .IN1(n1174), .IN3(n1172), .IN2(n1173), .IN4(n1171), .S0(N13), 
        .S1(n1424), .Q(n1175) );
  MUX41X1 U1401 ( .IN1(\mem[12][7] ), .IN3(\mem[14][7] ), .IN2(\mem[13][7] ), 
        .IN4(\mem[15][7] ), .S0(n1432), .S1(n1451), .Q(n1176) );
  MUX41X1 U1402 ( .IN1(\mem[8][7] ), .IN3(\mem[10][7] ), .IN2(\mem[9][7] ), 
        .IN4(\mem[11][7] ), .S0(n1432), .S1(n1451), .Q(n1177) );
  MUX41X1 U1403 ( .IN1(\mem[4][7] ), .IN3(\mem[6][7] ), .IN2(\mem[5][7] ), 
        .IN4(\mem[7][7] ), .S0(n1432), .S1(n1451), .Q(n1178) );
  MUX41X1 U1404 ( .IN1(\mem[0][7] ), .IN3(\mem[2][7] ), .IN2(\mem[1][7] ), 
        .IN4(\mem[3][7] ), .S0(n1432), .S1(n1451), .Q(n1179) );
  MUX41X1 U1405 ( .IN1(n1179), .IN3(n1177), .IN2(n1178), .IN4(n1176), .S0(N13), 
        .S1(n1424), .Q(n1180) );
  MUX21X1 U1406 ( .IN1(n1180), .IN2(n1175), .S(N14), .Q(rd_dataA[7]) );
  MUX41X1 U1407 ( .IN1(\mem[28][8] ), .IN3(\mem[30][8] ), .IN2(\mem[29][8] ), 
        .IN4(\mem[31][8] ), .S0(n1433), .S1(n1452), .Q(n1181) );
  MUX41X1 U1408 ( .IN1(\mem[24][8] ), .IN3(\mem[26][8] ), .IN2(\mem[25][8] ), 
        .IN4(\mem[27][8] ), .S0(n1433), .S1(n1452), .Q(n1182) );
  MUX41X1 U1409 ( .IN1(\mem[20][8] ), .IN3(\mem[22][8] ), .IN2(\mem[21][8] ), 
        .IN4(\mem[23][8] ), .S0(n1433), .S1(n1452), .Q(n1183) );
  MUX41X1 U1410 ( .IN1(\mem[16][8] ), .IN3(\mem[18][8] ), .IN2(\mem[17][8] ), 
        .IN4(\mem[19][8] ), .S0(n1433), .S1(n1452), .Q(n1184) );
  MUX41X1 U1411 ( .IN1(n1184), .IN3(n1182), .IN2(n1183), .IN4(n1181), .S0(N13), 
        .S1(n1424), .Q(n1185) );
  MUX41X1 U1412 ( .IN1(\mem[12][8] ), .IN3(\mem[14][8] ), .IN2(\mem[13][8] ), 
        .IN4(\mem[15][8] ), .S0(n1433), .S1(n1452), .Q(n1186) );
  MUX41X1 U1413 ( .IN1(\mem[8][8] ), .IN3(\mem[10][8] ), .IN2(\mem[9][8] ), 
        .IN4(\mem[11][8] ), .S0(n1433), .S1(n1452), .Q(n1187) );
  MUX41X1 U1414 ( .IN1(\mem[4][8] ), .IN3(\mem[6][8] ), .IN2(\mem[5][8] ), 
        .IN4(\mem[7][8] ), .S0(n1433), .S1(n1452), .Q(n1188) );
  MUX41X1 U1415 ( .IN1(\mem[0][8] ), .IN3(\mem[2][8] ), .IN2(\mem[1][8] ), 
        .IN4(\mem[3][8] ), .S0(n1433), .S1(n1452), .Q(n1189) );
  MUX41X1 U1416 ( .IN1(n1189), .IN3(n1187), .IN2(n1188), .IN4(n1186), .S0(N13), 
        .S1(n1424), .Q(n1190) );
  MUX21X1 U1417 ( .IN1(n1190), .IN2(n1185), .S(N14), .Q(rd_dataA[8]) );
  MUX41X1 U1418 ( .IN1(\mem[28][9] ), .IN3(\mem[30][9] ), .IN2(\mem[29][9] ), 
        .IN4(\mem[31][9] ), .S0(n1433), .S1(n1452), .Q(n1191) );
  MUX41X1 U1419 ( .IN1(\mem[24][9] ), .IN3(\mem[26][9] ), .IN2(\mem[25][9] ), 
        .IN4(\mem[27][9] ), .S0(n1433), .S1(n1452), .Q(n1192) );
  MUX41X1 U1420 ( .IN1(\mem[20][9] ), .IN3(\mem[22][9] ), .IN2(\mem[21][9] ), 
        .IN4(\mem[23][9] ), .S0(n1433), .S1(n1452), .Q(n1193) );
  MUX41X1 U1421 ( .IN1(\mem[16][9] ), .IN3(\mem[18][9] ), .IN2(\mem[17][9] ), 
        .IN4(\mem[19][9] ), .S0(n1433), .S1(n1452), .Q(n1194) );
  MUX41X1 U1422 ( .IN1(n1194), .IN3(n1192), .IN2(n1193), .IN4(n1191), .S0(N13), 
        .S1(n1424), .Q(n1195) );
  MUX41X1 U1423 ( .IN1(\mem[12][9] ), .IN3(\mem[14][9] ), .IN2(\mem[13][9] ), 
        .IN4(\mem[15][9] ), .S0(n1434), .S1(n1453), .Q(n1196) );
  MUX41X1 U1424 ( .IN1(\mem[8][9] ), .IN3(\mem[10][9] ), .IN2(\mem[9][9] ), 
        .IN4(\mem[11][9] ), .S0(n1434), .S1(n1453), .Q(n1197) );
  MUX41X1 U1425 ( .IN1(\mem[4][9] ), .IN3(\mem[6][9] ), .IN2(\mem[5][9] ), 
        .IN4(\mem[7][9] ), .S0(n1434), .S1(n1453), .Q(n1198) );
  MUX41X1 U1426 ( .IN1(\mem[0][9] ), .IN3(\mem[2][9] ), .IN2(\mem[1][9] ), 
        .IN4(\mem[3][9] ), .S0(n1434), .S1(n1453), .Q(n1199) );
  MUX41X1 U1427 ( .IN1(n1199), .IN3(n1197), .IN2(n1198), .IN4(n1196), .S0(N13), 
        .S1(n1424), .Q(n1200) );
  MUX21X1 U1428 ( .IN1(n1200), .IN2(n1195), .S(N14), .Q(rd_dataA[9]) );
  MUX41X1 U1429 ( .IN1(\mem[28][10] ), .IN3(\mem[30][10] ), .IN2(\mem[29][10] ), .IN4(\mem[31][10] ), .S0(n1434), .S1(n1453), .Q(n1201) );
  MUX41X1 U1430 ( .IN1(\mem[24][10] ), .IN3(\mem[26][10] ), .IN2(\mem[25][10] ), .IN4(\mem[27][10] ), .S0(n1434), .S1(n1453), .Q(n1202) );
  MUX41X1 U1431 ( .IN1(\mem[20][10] ), .IN3(\mem[22][10] ), .IN2(\mem[21][10] ), .IN4(\mem[23][10] ), .S0(n1434), .S1(n1453), .Q(n1203) );
  MUX41X1 U1432 ( .IN1(\mem[16][10] ), .IN3(\mem[18][10] ), .IN2(\mem[17][10] ), .IN4(\mem[19][10] ), .S0(n1434), .S1(n1453), .Q(n1204) );
  MUX41X1 U1433 ( .IN1(n1204), .IN3(n1202), .IN2(n1203), .IN4(n1201), .S0(N13), 
        .S1(n1424), .Q(n1205) );
  MUX41X1 U1434 ( .IN1(\mem[12][10] ), .IN3(\mem[14][10] ), .IN2(\mem[13][10] ), .IN4(\mem[15][10] ), .S0(n1434), .S1(n1453), .Q(n1206) );
  MUX41X1 U1435 ( .IN1(\mem[8][10] ), .IN3(\mem[10][10] ), .IN2(\mem[9][10] ), 
        .IN4(\mem[11][10] ), .S0(n1434), .S1(n1453), .Q(n1207) );
  MUX41X1 U1436 ( .IN1(\mem[4][10] ), .IN3(\mem[6][10] ), .IN2(\mem[5][10] ), 
        .IN4(\mem[7][10] ), .S0(n1434), .S1(n1453), .Q(n1208) );
  MUX41X1 U1437 ( .IN1(\mem[0][10] ), .IN3(\mem[2][10] ), .IN2(\mem[1][10] ), 
        .IN4(\mem[3][10] ), .S0(n1434), .S1(n1453), .Q(n1209) );
  MUX41X1 U1438 ( .IN1(n1209), .IN3(n1207), .IN2(n1208), .IN4(n1206), .S0(N13), 
        .S1(n1424), .Q(n1210) );
  MUX21X1 U1439 ( .IN1(n1210), .IN2(n1205), .S(N14), .Q(rd_dataA[10]) );
  MUX41X1 U1440 ( .IN1(\mem[28][11] ), .IN3(\mem[30][11] ), .IN2(\mem[29][11] ), .IN4(\mem[31][11] ), .S0(n1435), .S1(n1454), .Q(n1211) );
  MUX41X1 U1441 ( .IN1(\mem[24][11] ), .IN3(\mem[26][11] ), .IN2(\mem[25][11] ), .IN4(\mem[27][11] ), .S0(n1435), .S1(n1454), .Q(n1212) );
  MUX41X1 U1442 ( .IN1(\mem[20][11] ), .IN3(\mem[22][11] ), .IN2(\mem[21][11] ), .IN4(\mem[23][11] ), .S0(n1435), .S1(n1454), .Q(n1213) );
  MUX41X1 U1443 ( .IN1(\mem[16][11] ), .IN3(\mem[18][11] ), .IN2(\mem[17][11] ), .IN4(\mem[19][11] ), .S0(n1435), .S1(n1454), .Q(n1214) );
  MUX41X1 U1444 ( .IN1(n1214), .IN3(n1212), .IN2(n1213), .IN4(n1211), .S0(N13), 
        .S1(n1424), .Q(n1215) );
  MUX41X1 U1445 ( .IN1(\mem[12][11] ), .IN3(\mem[14][11] ), .IN2(\mem[13][11] ), .IN4(\mem[15][11] ), .S0(n1435), .S1(n1454), .Q(n1216) );
  MUX41X1 U1446 ( .IN1(\mem[8][11] ), .IN3(\mem[10][11] ), .IN2(\mem[9][11] ), 
        .IN4(\mem[11][11] ), .S0(n1435), .S1(n1454), .Q(n1217) );
  MUX41X1 U1447 ( .IN1(\mem[4][11] ), .IN3(\mem[6][11] ), .IN2(\mem[5][11] ), 
        .IN4(\mem[7][11] ), .S0(n1435), .S1(n1454), .Q(n1218) );
  MUX41X1 U1448 ( .IN1(\mem[0][11] ), .IN3(\mem[2][11] ), .IN2(\mem[1][11] ), 
        .IN4(\mem[3][11] ), .S0(n1435), .S1(n1454), .Q(n1219) );
  MUX41X1 U1449 ( .IN1(n1219), .IN3(n1217), .IN2(n1218), .IN4(n1216), .S0(N13), 
        .S1(n1424), .Q(n1220) );
  MUX21X1 U1450 ( .IN1(n1220), .IN2(n1215), .S(N14), .Q(rd_dataA[11]) );
  MUX41X1 U1451 ( .IN1(\mem[28][12] ), .IN3(\mem[30][12] ), .IN2(\mem[29][12] ), .IN4(\mem[31][12] ), .S0(n1435), .S1(n1454), .Q(n1221) );
  MUX41X1 U1452 ( .IN1(\mem[24][12] ), .IN3(\mem[26][12] ), .IN2(\mem[25][12] ), .IN4(\mem[27][12] ), .S0(n1435), .S1(n1454), .Q(n1222) );
  MUX41X1 U1453 ( .IN1(\mem[20][12] ), .IN3(\mem[22][12] ), .IN2(\mem[21][12] ), .IN4(\mem[23][12] ), .S0(n1435), .S1(n1454), .Q(n1223) );
  MUX41X1 U1454 ( .IN1(\mem[16][12] ), .IN3(\mem[18][12] ), .IN2(\mem[17][12] ), .IN4(\mem[19][12] ), .S0(n1435), .S1(n1454), .Q(n1224) );
  MUX41X1 U1455 ( .IN1(n1224), .IN3(n1222), .IN2(n1223), .IN4(n1221), .S0(N13), 
        .S1(N12), .Q(n1225) );
  MUX41X1 U1456 ( .IN1(\mem[12][12] ), .IN3(\mem[14][12] ), .IN2(\mem[13][12] ), .IN4(\mem[15][12] ), .S0(n1436), .S1(n1455), .Q(n1226) );
  MUX41X1 U1457 ( .IN1(\mem[8][12] ), .IN3(\mem[10][12] ), .IN2(\mem[9][12] ), 
        .IN4(\mem[11][12] ), .S0(n1436), .S1(n1455), .Q(n1227) );
  MUX41X1 U1458 ( .IN1(\mem[4][12] ), .IN3(\mem[6][12] ), .IN2(\mem[5][12] ), 
        .IN4(\mem[7][12] ), .S0(n1436), .S1(n1455), .Q(n1228) );
  MUX41X1 U1459 ( .IN1(\mem[0][12] ), .IN3(\mem[2][12] ), .IN2(\mem[1][12] ), 
        .IN4(\mem[3][12] ), .S0(n1436), .S1(n1455), .Q(n1229) );
  MUX41X1 U1460 ( .IN1(n1229), .IN3(n1227), .IN2(n1228), .IN4(n1226), .S0(N13), 
        .S1(N12), .Q(n1230) );
  MUX21X1 U1461 ( .IN1(n1230), .IN2(n1225), .S(N14), .Q(rd_dataA[12]) );
  MUX41X1 U1462 ( .IN1(\mem[28][13] ), .IN3(\mem[30][13] ), .IN2(\mem[29][13] ), .IN4(\mem[31][13] ), .S0(n1436), .S1(n1455), .Q(n1231) );
  MUX41X1 U1463 ( .IN1(\mem[24][13] ), .IN3(\mem[26][13] ), .IN2(\mem[25][13] ), .IN4(\mem[27][13] ), .S0(n1436), .S1(n1455), .Q(n1232) );
  MUX41X1 U1464 ( .IN1(\mem[20][13] ), .IN3(\mem[22][13] ), .IN2(\mem[21][13] ), .IN4(\mem[23][13] ), .S0(n1436), .S1(n1455), .Q(n1233) );
  MUX41X1 U1465 ( .IN1(\mem[16][13] ), .IN3(\mem[18][13] ), .IN2(\mem[17][13] ), .IN4(\mem[19][13] ), .S0(n1436), .S1(n1455), .Q(n1234) );
  MUX41X1 U1466 ( .IN1(n1234), .IN3(n1232), .IN2(n1233), .IN4(n1231), .S0(N13), 
        .S1(N12), .Q(n1235) );
  MUX41X1 U1467 ( .IN1(\mem[12][13] ), .IN3(\mem[14][13] ), .IN2(\mem[13][13] ), .IN4(\mem[15][13] ), .S0(n1436), .S1(n1455), .Q(n1236) );
  MUX41X1 U1468 ( .IN1(\mem[8][13] ), .IN3(\mem[10][13] ), .IN2(\mem[9][13] ), 
        .IN4(\mem[11][13] ), .S0(n1436), .S1(n1455), .Q(n1237) );
  MUX41X1 U1469 ( .IN1(\mem[4][13] ), .IN3(\mem[6][13] ), .IN2(\mem[5][13] ), 
        .IN4(\mem[7][13] ), .S0(n1436), .S1(n1455), .Q(n1238) );
  MUX41X1 U1470 ( .IN1(\mem[0][13] ), .IN3(\mem[2][13] ), .IN2(\mem[1][13] ), 
        .IN4(\mem[3][13] ), .S0(n1436), .S1(n1455), .Q(n1239) );
  MUX41X1 U1471 ( .IN1(n1239), .IN3(n1237), .IN2(n1238), .IN4(n1236), .S0(N13), 
        .S1(N12), .Q(n1240) );
  MUX21X1 U1472 ( .IN1(n1240), .IN2(n1235), .S(N14), .Q(rd_dataA[13]) );
  MUX41X1 U1473 ( .IN1(\mem[28][14] ), .IN3(\mem[30][14] ), .IN2(\mem[29][14] ), .IN4(\mem[31][14] ), .S0(N11), .S1(n1456), .Q(n1241) );
  MUX41X1 U1474 ( .IN1(\mem[24][14] ), .IN3(\mem[26][14] ), .IN2(\mem[25][14] ), .IN4(\mem[27][14] ), .S0(n1434), .S1(n1453), .Q(n1242) );
  MUX41X1 U1475 ( .IN1(\mem[20][14] ), .IN3(\mem[22][14] ), .IN2(\mem[21][14] ), .IN4(\mem[23][14] ), .S0(n1430), .S1(n1449), .Q(n1243) );
  MUX41X1 U1476 ( .IN1(\mem[16][14] ), .IN3(\mem[18][14] ), .IN2(\mem[17][14] ), .IN4(\mem[19][14] ), .S0(n1428), .S1(n1447), .Q(n1244) );
  MUX41X1 U1477 ( .IN1(n1244), .IN3(n1242), .IN2(n1243), .IN4(n1241), .S0(N13), 
        .S1(N12), .Q(n1245) );
  MUX41X1 U1478 ( .IN1(\mem[12][14] ), .IN3(\mem[14][14] ), .IN2(\mem[13][14] ), .IN4(\mem[15][14] ), .S0(N11), .S1(N10), .Q(n1246) );
  MUX41X1 U1479 ( .IN1(\mem[8][14] ), .IN3(\mem[10][14] ), .IN2(\mem[9][14] ), 
        .IN4(\mem[11][14] ), .S0(n1436), .S1(n1455), .Q(n1247) );
  MUX41X1 U1480 ( .IN1(\mem[4][14] ), .IN3(\mem[6][14] ), .IN2(\mem[5][14] ), 
        .IN4(\mem[7][14] ), .S0(n1433), .S1(n1452), .Q(n1248) );
  MUX41X1 U1481 ( .IN1(\mem[0][14] ), .IN3(\mem[2][14] ), .IN2(\mem[1][14] ), 
        .IN4(\mem[3][14] ), .S0(n1432), .S1(n1451), .Q(n1249) );
  MUX41X1 U1482 ( .IN1(n1249), .IN3(n1247), .IN2(n1248), .IN4(n1246), .S0(N13), 
        .S1(N12), .Q(n1250) );
  MUX21X1 U1483 ( .IN1(n1250), .IN2(n1245), .S(N14), .Q(rd_dataA[14]) );
  MUX41X1 U1484 ( .IN1(\mem[28][15] ), .IN3(\mem[30][15] ), .IN2(\mem[29][15] ), .IN4(\mem[31][15] ), .S0(N11), .S1(N10), .Q(n1251) );
  MUX41X1 U1485 ( .IN1(\mem[24][15] ), .IN3(\mem[26][15] ), .IN2(\mem[25][15] ), .IN4(\mem[27][15] ), .S0(n1435), .S1(n1454), .Q(n1252) );
  MUX41X1 U1486 ( .IN1(\mem[20][15] ), .IN3(\mem[22][15] ), .IN2(\mem[21][15] ), .IN4(\mem[23][15] ), .S0(n1431), .S1(n1450), .Q(n1253) );
  MUX41X1 U1487 ( .IN1(\mem[16][15] ), .IN3(\mem[18][15] ), .IN2(\mem[17][15] ), .IN4(\mem[19][15] ), .S0(n1429), .S1(n1448), .Q(n1254) );
  MUX41X1 U1488 ( .IN1(n1254), .IN3(n1252), .IN2(n1253), .IN4(n1251), .S0(N13), 
        .S1(N12), .Q(n1255) );
  MUX41X1 U1489 ( .IN1(\mem[12][15] ), .IN3(\mem[14][15] ), .IN2(\mem[13][15] ), .IN4(\mem[15][15] ), .S0(n1438), .S1(n1456), .Q(n1256) );
  MUX41X1 U1490 ( .IN1(\mem[8][15] ), .IN3(\mem[10][15] ), .IN2(\mem[9][15] ), 
        .IN4(\mem[11][15] ), .S0(n1435), .S1(n1456), .Q(n1257) );
  MUX41X1 U1491 ( .IN1(\mem[4][15] ), .IN3(\mem[6][15] ), .IN2(\mem[5][15] ), 
        .IN4(\mem[7][15] ), .S0(n1432), .S1(n1456), .Q(n1258) );
  MUX41X1 U1492 ( .IN1(\mem[0][15] ), .IN3(\mem[2][15] ), .IN2(\mem[1][15] ), 
        .IN4(\mem[3][15] ), .S0(n1430), .S1(n1456), .Q(n1259) );
  MUX41X1 U1493 ( .IN1(n1259), .IN3(n1257), .IN2(n1258), .IN4(n1256), .S0(N13), 
        .S1(N12), .Q(n1260) );
  MUX21X1 U1494 ( .IN1(n1260), .IN2(n1255), .S(N14), .Q(rd_dataA[15]) );
  MUX41X1 U1495 ( .IN1(\mem[28][16] ), .IN3(\mem[30][16] ), .IN2(\mem[29][16] ), .IN4(\mem[31][16] ), .S0(N11), .S1(n1456), .Q(n1261) );
  MUX41X1 U1496 ( .IN1(\mem[24][16] ), .IN3(\mem[26][16] ), .IN2(\mem[25][16] ), .IN4(\mem[27][16] ), .S0(n1434), .S1(n1456), .Q(n1262) );
  MUX41X1 U1497 ( .IN1(\mem[20][16] ), .IN3(\mem[22][16] ), .IN2(\mem[21][16] ), .IN4(\mem[23][16] ), .S0(n1429), .S1(n1456), .Q(n1263) );
  MUX41X1 U1498 ( .IN1(\mem[16][16] ), .IN3(\mem[18][16] ), .IN2(\mem[17][16] ), .IN4(\mem[19][16] ), .S0(n1428), .S1(n1456), .Q(n1264) );
  MUX41X1 U1499 ( .IN1(n1264), .IN3(n1262), .IN2(n1263), .IN4(n1261), .S0(N13), 
        .S1(n1424), .Q(n1265) );
  MUX41X1 U1500 ( .IN1(\mem[12][16] ), .IN3(\mem[14][16] ), .IN2(\mem[13][16] ), .IN4(\mem[15][16] ), .S0(n1439), .S1(n1456), .Q(n1266) );
  MUX41X1 U1501 ( .IN1(\mem[8][16] ), .IN3(\mem[10][16] ), .IN2(\mem[9][16] ), 
        .IN4(\mem[11][16] ), .S0(n1436), .S1(n1456), .Q(n1267) );
  MUX41X1 U1502 ( .IN1(\mem[4][16] ), .IN3(\mem[6][16] ), .IN2(\mem[5][16] ), 
        .IN4(\mem[7][16] ), .S0(n1433), .S1(n1456), .Q(n1268) );
  MUX41X1 U1503 ( .IN1(\mem[0][16] ), .IN3(\mem[2][16] ), .IN2(\mem[1][16] ), 
        .IN4(\mem[3][16] ), .S0(n1431), .S1(n1456), .Q(n1269) );
  MUX41X1 U1504 ( .IN1(n1269), .IN3(n1267), .IN2(n1268), .IN4(n1266), .S0(N13), 
        .S1(N12), .Q(n1270) );
  MUX21X1 U1505 ( .IN1(n1270), .IN2(n1265), .S(N14), .Q(rd_dataA[16]) );
  MUX41X1 U1506 ( .IN1(\mem[28][17] ), .IN3(\mem[30][17] ), .IN2(\mem[29][17] ), .IN4(\mem[31][17] ), .S0(n1437), .S1(n1457), .Q(n1271) );
  MUX41X1 U1507 ( .IN1(\mem[24][17] ), .IN3(\mem[26][17] ), .IN2(\mem[25][17] ), .IN4(\mem[27][17] ), .S0(n1437), .S1(n1457), .Q(n1272) );
  MUX41X1 U1508 ( .IN1(\mem[20][17] ), .IN3(\mem[22][17] ), .IN2(\mem[21][17] ), .IN4(\mem[23][17] ), .S0(n1437), .S1(n1457), .Q(n1273) );
  MUX41X1 U1509 ( .IN1(\mem[16][17] ), .IN3(\mem[18][17] ), .IN2(\mem[17][17] ), .IN4(\mem[19][17] ), .S0(n1437), .S1(n1457), .Q(n1274) );
  MUX41X1 U1510 ( .IN1(n1274), .IN3(n1272), .IN2(n1273), .IN4(n1271), .S0(N13), 
        .S1(n1425), .Q(n1275) );
  MUX41X1 U1511 ( .IN1(\mem[12][17] ), .IN3(\mem[14][17] ), .IN2(\mem[13][17] ), .IN4(\mem[15][17] ), .S0(n1437), .S1(n1457), .Q(n1276) );
  MUX41X1 U1512 ( .IN1(\mem[8][17] ), .IN3(\mem[10][17] ), .IN2(\mem[9][17] ), 
        .IN4(\mem[11][17] ), .S0(n1437), .S1(n1457), .Q(n1277) );
  MUX41X1 U1513 ( .IN1(\mem[4][17] ), .IN3(\mem[6][17] ), .IN2(\mem[5][17] ), 
        .IN4(\mem[7][17] ), .S0(n1437), .S1(n1457), .Q(n1278) );
  MUX41X1 U1514 ( .IN1(\mem[0][17] ), .IN3(\mem[2][17] ), .IN2(\mem[1][17] ), 
        .IN4(\mem[3][17] ), .S0(n1437), .S1(n1457), .Q(n1279) );
  MUX41X1 U1515 ( .IN1(n1279), .IN3(n1277), .IN2(n1278), .IN4(n1276), .S0(N13), 
        .S1(N12), .Q(n1280) );
  MUX21X1 U1516 ( .IN1(n1280), .IN2(n1275), .S(N14), .Q(rd_dataA[17]) );
  MUX41X1 U1517 ( .IN1(\mem[28][18] ), .IN3(\mem[30][18] ), .IN2(\mem[29][18] ), .IN4(\mem[31][18] ), .S0(n1437), .S1(n1457), .Q(n1281) );
  MUX41X1 U1518 ( .IN1(\mem[24][18] ), .IN3(\mem[26][18] ), .IN2(\mem[25][18] ), .IN4(\mem[27][18] ), .S0(n1437), .S1(n1457), .Q(n1282) );
  MUX41X1 U1519 ( .IN1(\mem[20][18] ), .IN3(\mem[22][18] ), .IN2(\mem[21][18] ), .IN4(\mem[23][18] ), .S0(n1437), .S1(n1457), .Q(n1283) );
  MUX41X1 U1520 ( .IN1(\mem[16][18] ), .IN3(\mem[18][18] ), .IN2(\mem[17][18] ), .IN4(\mem[19][18] ), .S0(n1437), .S1(n1457), .Q(n1284) );
  MUX41X1 U1521 ( .IN1(n1284), .IN3(n1282), .IN2(n1283), .IN4(n1281), .S0(N13), 
        .S1(n1423), .Q(n1285) );
  MUX41X1 U1522 ( .IN1(\mem[12][18] ), .IN3(\mem[14][18] ), .IN2(\mem[13][18] ), .IN4(\mem[15][18] ), .S0(n1438), .S1(n1458), .Q(n1286) );
  MUX41X1 U1523 ( .IN1(\mem[8][18] ), .IN3(\mem[10][18] ), .IN2(\mem[9][18] ), 
        .IN4(\mem[11][18] ), .S0(n1438), .S1(n1458), .Q(n1287) );
  MUX41X1 U1524 ( .IN1(\mem[4][18] ), .IN3(\mem[6][18] ), .IN2(\mem[5][18] ), 
        .IN4(\mem[7][18] ), .S0(n1438), .S1(n1458), .Q(n1288) );
  MUX41X1 U1525 ( .IN1(\mem[0][18] ), .IN3(\mem[2][18] ), .IN2(\mem[1][18] ), 
        .IN4(\mem[3][18] ), .S0(n1438), .S1(n1458), .Q(n1289) );
  MUX41X1 U1526 ( .IN1(n1289), .IN3(n1287), .IN2(n1288), .IN4(n1286), .S0(N13), 
        .S1(n1423), .Q(n1290) );
  MUX21X1 U1527 ( .IN1(n1290), .IN2(n1285), .S(N14), .Q(rd_dataA[18]) );
  MUX41X1 U1528 ( .IN1(\mem[28][19] ), .IN3(\mem[30][19] ), .IN2(\mem[29][19] ), .IN4(\mem[31][19] ), .S0(n1438), .S1(n1458), .Q(n1291) );
  MUX41X1 U1529 ( .IN1(\mem[24][19] ), .IN3(\mem[26][19] ), .IN2(\mem[25][19] ), .IN4(\mem[27][19] ), .S0(n1438), .S1(n1458), .Q(n1292) );
  MUX41X1 U1530 ( .IN1(\mem[20][19] ), .IN3(\mem[22][19] ), .IN2(\mem[21][19] ), .IN4(\mem[23][19] ), .S0(n1438), .S1(n1458), .Q(n1293) );
  MUX41X1 U1531 ( .IN1(\mem[16][19] ), .IN3(\mem[18][19] ), .IN2(\mem[17][19] ), .IN4(\mem[19][19] ), .S0(n1438), .S1(n1458), .Q(n1294) );
  MUX41X1 U1532 ( .IN1(n1294), .IN3(n1292), .IN2(n1293), .IN4(n1291), .S0(N13), 
        .S1(n1423), .Q(n1295) );
  MUX41X1 U1533 ( .IN1(\mem[12][19] ), .IN3(\mem[14][19] ), .IN2(\mem[13][19] ), .IN4(\mem[15][19] ), .S0(n1438), .S1(n1458), .Q(n1296) );
  MUX41X1 U1534 ( .IN1(\mem[8][19] ), .IN3(\mem[10][19] ), .IN2(\mem[9][19] ), 
        .IN4(\mem[11][19] ), .S0(n1438), .S1(n1458), .Q(n1297) );
  MUX41X1 U1535 ( .IN1(\mem[4][19] ), .IN3(\mem[6][19] ), .IN2(\mem[5][19] ), 
        .IN4(\mem[7][19] ), .S0(n1438), .S1(n1458), .Q(n1298) );
  MUX41X1 U1536 ( .IN1(\mem[0][19] ), .IN3(\mem[2][19] ), .IN2(\mem[1][19] ), 
        .IN4(\mem[3][19] ), .S0(n1438), .S1(n1458), .Q(n1299) );
  MUX41X1 U1537 ( .IN1(n1299), .IN3(n1297), .IN2(n1298), .IN4(n1296), .S0(N13), 
        .S1(n1423), .Q(n1300) );
  MUX21X1 U1538 ( .IN1(n1300), .IN2(n1295), .S(N14), .Q(rd_dataA[19]) );
  MUX41X1 U1539 ( .IN1(\mem[28][20] ), .IN3(\mem[30][20] ), .IN2(\mem[29][20] ), .IN4(\mem[31][20] ), .S0(n1439), .S1(n1459), .Q(n1301) );
  MUX41X1 U1540 ( .IN1(\mem[24][20] ), .IN3(\mem[26][20] ), .IN2(\mem[25][20] ), .IN4(\mem[27][20] ), .S0(n1439), .S1(n1459), .Q(n1302) );
  MUX41X1 U1541 ( .IN1(\mem[20][20] ), .IN3(\mem[22][20] ), .IN2(\mem[21][20] ), .IN4(\mem[23][20] ), .S0(n1439), .S1(n1459), .Q(n1303) );
  MUX41X1 U1542 ( .IN1(\mem[16][20] ), .IN3(\mem[18][20] ), .IN2(\mem[17][20] ), .IN4(\mem[19][20] ), .S0(n1439), .S1(n1459), .Q(n1304) );
  MUX41X1 U1543 ( .IN1(n1304), .IN3(n1302), .IN2(n1303), .IN4(n1301), .S0(N13), 
        .S1(n1423), .Q(n1305) );
  MUX41X1 U1544 ( .IN1(\mem[12][20] ), .IN3(\mem[14][20] ), .IN2(\mem[13][20] ), .IN4(\mem[15][20] ), .S0(n1439), .S1(n1459), .Q(n1306) );
  MUX41X1 U1545 ( .IN1(\mem[8][20] ), .IN3(\mem[10][20] ), .IN2(\mem[9][20] ), 
        .IN4(\mem[11][20] ), .S0(n1439), .S1(n1459), .Q(n1307) );
  MUX41X1 U1546 ( .IN1(\mem[4][20] ), .IN3(\mem[6][20] ), .IN2(\mem[5][20] ), 
        .IN4(\mem[7][20] ), .S0(n1439), .S1(n1459), .Q(n1308) );
  MUX41X1 U1547 ( .IN1(\mem[0][20] ), .IN3(\mem[2][20] ), .IN2(\mem[1][20] ), 
        .IN4(\mem[3][20] ), .S0(n1439), .S1(n1459), .Q(n1309) );
  MUX41X1 U1548 ( .IN1(n1309), .IN3(n1307), .IN2(n1308), .IN4(n1306), .S0(N13), 
        .S1(n1423), .Q(n1310) );
  MUX21X1 U1549 ( .IN1(n1310), .IN2(n1305), .S(N14), .Q(rd_dataA[20]) );
  MUX41X1 U1550 ( .IN1(\mem[28][21] ), .IN3(\mem[30][21] ), .IN2(\mem[29][21] ), .IN4(\mem[31][21] ), .S0(n1439), .S1(n1459), .Q(n1311) );
  MUX41X1 U1551 ( .IN1(\mem[24][21] ), .IN3(\mem[26][21] ), .IN2(\mem[25][21] ), .IN4(\mem[27][21] ), .S0(n1439), .S1(n1459), .Q(n1312) );
  MUX41X1 U1552 ( .IN1(\mem[20][21] ), .IN3(\mem[22][21] ), .IN2(\mem[21][21] ), .IN4(\mem[23][21] ), .S0(n1439), .S1(n1459), .Q(n1313) );
  MUX41X1 U1553 ( .IN1(\mem[16][21] ), .IN3(\mem[18][21] ), .IN2(\mem[17][21] ), .IN4(\mem[19][21] ), .S0(n1439), .S1(n1459), .Q(n1314) );
  MUX41X1 U1554 ( .IN1(n1314), .IN3(n1312), .IN2(n1313), .IN4(n1311), .S0(N13), 
        .S1(n1423), .Q(n1315) );
  MUX41X1 U1555 ( .IN1(\mem[12][21] ), .IN3(\mem[14][21] ), .IN2(\mem[13][21] ), .IN4(\mem[15][21] ), .S0(n1440), .S1(n1460), .Q(n1316) );
  MUX41X1 U1556 ( .IN1(\mem[8][21] ), .IN3(\mem[10][21] ), .IN2(\mem[9][21] ), 
        .IN4(\mem[11][21] ), .S0(n1440), .S1(n1460), .Q(n1317) );
  MUX41X1 U1557 ( .IN1(\mem[4][21] ), .IN3(\mem[6][21] ), .IN2(\mem[5][21] ), 
        .IN4(\mem[7][21] ), .S0(n1440), .S1(n1460), .Q(n1318) );
  MUX41X1 U1558 ( .IN1(\mem[0][21] ), .IN3(\mem[2][21] ), .IN2(\mem[1][21] ), 
        .IN4(\mem[3][21] ), .S0(n1440), .S1(n1460), .Q(n1319) );
  MUX41X1 U1559 ( .IN1(n1319), .IN3(n1317), .IN2(n1318), .IN4(n1316), .S0(N13), 
        .S1(n1423), .Q(n1320) );
  MUX21X1 U1560 ( .IN1(n1320), .IN2(n1315), .S(N14), .Q(rd_dataA[21]) );
  MUX41X1 U1561 ( .IN1(\mem[28][22] ), .IN3(\mem[30][22] ), .IN2(\mem[29][22] ), .IN4(\mem[31][22] ), .S0(n1440), .S1(n1460), .Q(n1321) );
  MUX41X1 U1562 ( .IN1(\mem[24][22] ), .IN3(\mem[26][22] ), .IN2(\mem[25][22] ), .IN4(\mem[27][22] ), .S0(n1440), .S1(n1460), .Q(n1322) );
  MUX41X1 U1563 ( .IN1(\mem[20][22] ), .IN3(\mem[22][22] ), .IN2(\mem[21][22] ), .IN4(\mem[23][22] ), .S0(n1440), .S1(n1460), .Q(n1323) );
  MUX41X1 U1564 ( .IN1(\mem[16][22] ), .IN3(\mem[18][22] ), .IN2(\mem[17][22] ), .IN4(\mem[19][22] ), .S0(n1440), .S1(n1460), .Q(n1324) );
  MUX41X1 U1565 ( .IN1(n1324), .IN3(n1322), .IN2(n1323), .IN4(n1321), .S0(N13), 
        .S1(n1423), .Q(n1325) );
  MUX41X1 U1566 ( .IN1(\mem[12][22] ), .IN3(\mem[14][22] ), .IN2(\mem[13][22] ), .IN4(\mem[15][22] ), .S0(n1440), .S1(n1460), .Q(n1326) );
  MUX41X1 U1567 ( .IN1(\mem[8][22] ), .IN3(\mem[10][22] ), .IN2(\mem[9][22] ), 
        .IN4(\mem[11][22] ), .S0(n1440), .S1(n1460), .Q(n1327) );
  MUX41X1 U1568 ( .IN1(\mem[4][22] ), .IN3(\mem[6][22] ), .IN2(\mem[5][22] ), 
        .IN4(\mem[7][22] ), .S0(n1440), .S1(n1460), .Q(n1328) );
  MUX41X1 U1569 ( .IN1(\mem[0][22] ), .IN3(\mem[2][22] ), .IN2(\mem[1][22] ), 
        .IN4(\mem[3][22] ), .S0(n1440), .S1(n1460), .Q(n1329) );
  MUX41X1 U1570 ( .IN1(n1329), .IN3(n1327), .IN2(n1328), .IN4(n1326), .S0(N13), 
        .S1(n1423), .Q(n1330) );
  MUX21X1 U1571 ( .IN1(n1330), .IN2(n1325), .S(N14), .Q(rd_dataA[22]) );
  MUX41X1 U1572 ( .IN1(\mem[28][23] ), .IN3(\mem[30][23] ), .IN2(\mem[29][23] ), .IN4(\mem[31][23] ), .S0(n1441), .S1(n1461), .Q(n1331) );
  MUX41X1 U1573 ( .IN1(\mem[24][23] ), .IN3(\mem[26][23] ), .IN2(\mem[25][23] ), .IN4(\mem[27][23] ), .S0(n1441), .S1(n1461), .Q(n1332) );
  MUX41X1 U1574 ( .IN1(\mem[20][23] ), .IN3(\mem[22][23] ), .IN2(\mem[21][23] ), .IN4(\mem[23][23] ), .S0(n1441), .S1(n1461), .Q(n1333) );
  MUX41X1 U1575 ( .IN1(\mem[16][23] ), .IN3(\mem[18][23] ), .IN2(\mem[17][23] ), .IN4(\mem[19][23] ), .S0(n1441), .S1(n1461), .Q(n1334) );
  MUX41X1 U1576 ( .IN1(n1334), .IN3(n1332), .IN2(n1333), .IN4(n1331), .S0(N13), 
        .S1(n1423), .Q(n1335) );
  MUX41X1 U1577 ( .IN1(\mem[12][23] ), .IN3(\mem[14][23] ), .IN2(\mem[13][23] ), .IN4(\mem[15][23] ), .S0(n1441), .S1(n1461), .Q(n1336) );
  MUX41X1 U1578 ( .IN1(\mem[8][23] ), .IN3(\mem[10][23] ), .IN2(\mem[9][23] ), 
        .IN4(\mem[11][23] ), .S0(n1441), .S1(n1461), .Q(n1337) );
  MUX41X1 U1579 ( .IN1(\mem[4][23] ), .IN3(\mem[6][23] ), .IN2(\mem[5][23] ), 
        .IN4(\mem[7][23] ), .S0(n1441), .S1(n1461), .Q(n1338) );
  MUX41X1 U1580 ( .IN1(\mem[0][23] ), .IN3(\mem[2][23] ), .IN2(\mem[1][23] ), 
        .IN4(\mem[3][23] ), .S0(n1441), .S1(n1461), .Q(n1339) );
  MUX41X1 U1581 ( .IN1(n1339), .IN3(n1337), .IN2(n1338), .IN4(n1336), .S0(N13), 
        .S1(n1423), .Q(n1340) );
  MUX21X1 U1582 ( .IN1(n1340), .IN2(n1335), .S(N14), .Q(rd_dataA[23]) );
  MUX41X1 U1583 ( .IN1(\mem[28][24] ), .IN3(\mem[30][24] ), .IN2(\mem[29][24] ), .IN4(\mem[31][24] ), .S0(n1441), .S1(n1461), .Q(n1341) );
  MUX41X1 U1584 ( .IN1(\mem[24][24] ), .IN3(\mem[26][24] ), .IN2(\mem[25][24] ), .IN4(\mem[27][24] ), .S0(n1441), .S1(n1461), .Q(n1342) );
  MUX41X1 U1585 ( .IN1(\mem[20][24] ), .IN3(\mem[22][24] ), .IN2(\mem[21][24] ), .IN4(\mem[23][24] ), .S0(n1441), .S1(n1461), .Q(n1343) );
  MUX41X1 U1586 ( .IN1(\mem[16][24] ), .IN3(\mem[18][24] ), .IN2(\mem[17][24] ), .IN4(\mem[19][24] ), .S0(n1441), .S1(n1461), .Q(n1344) );
  MUX41X1 U1587 ( .IN1(n1344), .IN3(n1342), .IN2(n1343), .IN4(n1341), .S0(N13), 
        .S1(n1422), .Q(n1345) );
  MUX41X1 U1588 ( .IN1(\mem[12][24] ), .IN3(\mem[14][24] ), .IN2(\mem[13][24] ), .IN4(\mem[15][24] ), .S0(n1442), .S1(n1462), .Q(n1346) );
  MUX41X1 U1589 ( .IN1(\mem[8][24] ), .IN3(\mem[10][24] ), .IN2(\mem[9][24] ), 
        .IN4(\mem[11][24] ), .S0(n1442), .S1(n1462), .Q(n1347) );
  MUX41X1 U1590 ( .IN1(\mem[4][24] ), .IN3(\mem[6][24] ), .IN2(\mem[5][24] ), 
        .IN4(\mem[7][24] ), .S0(n1442), .S1(n1462), .Q(n1348) );
  MUX41X1 U1591 ( .IN1(\mem[0][24] ), .IN3(\mem[2][24] ), .IN2(\mem[1][24] ), 
        .IN4(\mem[3][24] ), .S0(n1442), .S1(n1462), .Q(n1349) );
  MUX41X1 U1592 ( .IN1(n1349), .IN3(n1347), .IN2(n1348), .IN4(n1346), .S0(N13), 
        .S1(n1422), .Q(n1350) );
  MUX21X1 U1593 ( .IN1(n1350), .IN2(n1345), .S(N14), .Q(rd_dataA[24]) );
  MUX41X1 U1594 ( .IN1(\mem[28][25] ), .IN3(\mem[30][25] ), .IN2(\mem[29][25] ), .IN4(\mem[31][25] ), .S0(n1442), .S1(n1462), .Q(n1351) );
  MUX41X1 U1595 ( .IN1(\mem[24][25] ), .IN3(\mem[26][25] ), .IN2(\mem[25][25] ), .IN4(\mem[27][25] ), .S0(n1442), .S1(n1462), .Q(n1352) );
  MUX41X1 U1596 ( .IN1(\mem[20][25] ), .IN3(\mem[22][25] ), .IN2(\mem[21][25] ), .IN4(\mem[23][25] ), .S0(n1442), .S1(n1462), .Q(n1353) );
  MUX41X1 U1597 ( .IN1(\mem[16][25] ), .IN3(\mem[18][25] ), .IN2(\mem[17][25] ), .IN4(\mem[19][25] ), .S0(n1442), .S1(n1462), .Q(n1354) );
  MUX41X1 U1598 ( .IN1(n1354), .IN3(n1352), .IN2(n1353), .IN4(n1351), .S0(N13), 
        .S1(n1422), .Q(n1355) );
  MUX41X1 U1599 ( .IN1(\mem[12][25] ), .IN3(\mem[14][25] ), .IN2(\mem[13][25] ), .IN4(\mem[15][25] ), .S0(n1442), .S1(n1462), .Q(n1356) );
  MUX41X1 U1600 ( .IN1(\mem[8][25] ), .IN3(\mem[10][25] ), .IN2(\mem[9][25] ), 
        .IN4(\mem[11][25] ), .S0(n1442), .S1(n1462), .Q(n1357) );
  MUX41X1 U1601 ( .IN1(\mem[4][25] ), .IN3(\mem[6][25] ), .IN2(\mem[5][25] ), 
        .IN4(\mem[7][25] ), .S0(n1442), .S1(n1462), .Q(n1358) );
  MUX41X1 U1602 ( .IN1(\mem[0][25] ), .IN3(\mem[2][25] ), .IN2(\mem[1][25] ), 
        .IN4(\mem[3][25] ), .S0(n1442), .S1(n1462), .Q(n1359) );
  MUX41X1 U1603 ( .IN1(n1359), .IN3(n1357), .IN2(n1358), .IN4(n1356), .S0(N13), 
        .S1(n1422), .Q(n1360) );
  MUX21X1 U1604 ( .IN1(n1360), .IN2(n1355), .S(N14), .Q(rd_dataA[25]) );
  MUX41X1 U1605 ( .IN1(\mem[28][26] ), .IN3(\mem[30][26] ), .IN2(\mem[29][26] ), .IN4(\mem[31][26] ), .S0(n1443), .S1(n1463), .Q(n1361) );
  MUX41X1 U1606 ( .IN1(\mem[24][26] ), .IN3(\mem[26][26] ), .IN2(\mem[25][26] ), .IN4(\mem[27][26] ), .S0(n1443), .S1(n1463), .Q(n1362) );
  MUX41X1 U1607 ( .IN1(\mem[20][26] ), .IN3(\mem[22][26] ), .IN2(\mem[21][26] ), .IN4(\mem[23][26] ), .S0(n1443), .S1(n1463), .Q(n1363) );
  MUX41X1 U1608 ( .IN1(\mem[16][26] ), .IN3(\mem[18][26] ), .IN2(\mem[17][26] ), .IN4(\mem[19][26] ), .S0(n1443), .S1(n1463), .Q(n1364) );
  MUX41X1 U1609 ( .IN1(n1364), .IN3(n1362), .IN2(n1363), .IN4(n1361), .S0(N13), 
        .S1(n1422), .Q(n1365) );
  MUX41X1 U1610 ( .IN1(\mem[12][26] ), .IN3(\mem[14][26] ), .IN2(\mem[13][26] ), .IN4(\mem[15][26] ), .S0(n1443), .S1(n1463), .Q(n1366) );
  MUX41X1 U1611 ( .IN1(\mem[8][26] ), .IN3(\mem[10][26] ), .IN2(\mem[9][26] ), 
        .IN4(\mem[11][26] ), .S0(n1443), .S1(n1463), .Q(n1367) );
  MUX41X1 U1612 ( .IN1(\mem[4][26] ), .IN3(\mem[6][26] ), .IN2(\mem[5][26] ), 
        .IN4(\mem[7][26] ), .S0(n1443), .S1(n1463), .Q(n1368) );
  MUX41X1 U1613 ( .IN1(\mem[0][26] ), .IN3(\mem[2][26] ), .IN2(\mem[1][26] ), 
        .IN4(\mem[3][26] ), .S0(n1443), .S1(n1463), .Q(n1369) );
  MUX41X1 U1614 ( .IN1(n1369), .IN3(n1367), .IN2(n1368), .IN4(n1366), .S0(N13), 
        .S1(n1422), .Q(n1370) );
  MUX21X1 U1615 ( .IN1(n1370), .IN2(n1365), .S(N14), .Q(rd_dataA[26]) );
  MUX41X1 U1616 ( .IN1(\mem[28][27] ), .IN3(\mem[30][27] ), .IN2(\mem[29][27] ), .IN4(\mem[31][27] ), .S0(n1443), .S1(n1463), .Q(n1371) );
  MUX41X1 U1617 ( .IN1(\mem[24][27] ), .IN3(\mem[26][27] ), .IN2(\mem[25][27] ), .IN4(\mem[27][27] ), .S0(n1443), .S1(n1463), .Q(n1372) );
  MUX41X1 U1618 ( .IN1(\mem[20][27] ), .IN3(\mem[22][27] ), .IN2(\mem[21][27] ), .IN4(\mem[23][27] ), .S0(n1443), .S1(n1463), .Q(n1373) );
  MUX41X1 U1619 ( .IN1(\mem[16][27] ), .IN3(\mem[18][27] ), .IN2(\mem[17][27] ), .IN4(\mem[19][27] ), .S0(n1443), .S1(n1463), .Q(n1374) );
  MUX41X1 U1620 ( .IN1(n1374), .IN3(n1372), .IN2(n1373), .IN4(n1371), .S0(N13), 
        .S1(n1422), .Q(n1375) );
  MUX41X1 U1621 ( .IN1(\mem[12][27] ), .IN3(\mem[14][27] ), .IN2(\mem[13][27] ), .IN4(\mem[15][27] ), .S0(n1444), .S1(n1464), .Q(n1376) );
  MUX41X1 U1622 ( .IN1(\mem[8][27] ), .IN3(\mem[10][27] ), .IN2(\mem[9][27] ), 
        .IN4(\mem[11][27] ), .S0(n1444), .S1(n1464), .Q(n1377) );
  MUX41X1 U1623 ( .IN1(\mem[4][27] ), .IN3(\mem[6][27] ), .IN2(\mem[5][27] ), 
        .IN4(\mem[7][27] ), .S0(n1444), .S1(n1464), .Q(n1378) );
  MUX41X1 U1624 ( .IN1(\mem[0][27] ), .IN3(\mem[2][27] ), .IN2(\mem[1][27] ), 
        .IN4(\mem[3][27] ), .S0(n1444), .S1(n1464), .Q(n1379) );
  MUX41X1 U1625 ( .IN1(n1379), .IN3(n1377), .IN2(n1378), .IN4(n1376), .S0(N13), 
        .S1(n1422), .Q(n1380) );
  MUX21X1 U1626 ( .IN1(n1380), .IN2(n1375), .S(N14), .Q(rd_dataA[27]) );
  MUX41X1 U1627 ( .IN1(\mem[28][28] ), .IN3(\mem[30][28] ), .IN2(\mem[29][28] ), .IN4(\mem[31][28] ), .S0(n1444), .S1(n1464), .Q(n1381) );
  MUX41X1 U1628 ( .IN1(\mem[24][28] ), .IN3(\mem[26][28] ), .IN2(\mem[25][28] ), .IN4(\mem[27][28] ), .S0(n1444), .S1(n1464), .Q(n1382) );
  MUX41X1 U1629 ( .IN1(\mem[20][28] ), .IN3(\mem[22][28] ), .IN2(\mem[21][28] ), .IN4(\mem[23][28] ), .S0(n1444), .S1(n1464), .Q(n1383) );
  MUX41X1 U1630 ( .IN1(\mem[16][28] ), .IN3(\mem[18][28] ), .IN2(\mem[17][28] ), .IN4(\mem[19][28] ), .S0(n1444), .S1(n1464), .Q(n1384) );
  MUX41X1 U1631 ( .IN1(n1384), .IN3(n1382), .IN2(n1383), .IN4(n1381), .S0(N13), 
        .S1(n1422), .Q(n1385) );
  MUX41X1 U1632 ( .IN1(\mem[12][28] ), .IN3(\mem[14][28] ), .IN2(\mem[13][28] ), .IN4(\mem[15][28] ), .S0(n1444), .S1(n1464), .Q(n1386) );
  MUX41X1 U1633 ( .IN1(\mem[8][28] ), .IN3(\mem[10][28] ), .IN2(\mem[9][28] ), 
        .IN4(\mem[11][28] ), .S0(n1444), .S1(n1464), .Q(n1387) );
  MUX41X1 U1634 ( .IN1(\mem[4][28] ), .IN3(\mem[6][28] ), .IN2(\mem[5][28] ), 
        .IN4(\mem[7][28] ), .S0(n1444), .S1(n1464), .Q(n1388) );
  MUX41X1 U1635 ( .IN1(\mem[0][28] ), .IN3(\mem[2][28] ), .IN2(\mem[1][28] ), 
        .IN4(\mem[3][28] ), .S0(n1444), .S1(n1464), .Q(n1389) );
  MUX41X1 U1636 ( .IN1(n1389), .IN3(n1387), .IN2(n1388), .IN4(n1386), .S0(N13), 
        .S1(n1422), .Q(n1390) );
  MUX21X1 U1637 ( .IN1(n1390), .IN2(n1385), .S(N14), .Q(rd_dataA[28]) );
  MUX41X1 U1638 ( .IN1(\mem[28][29] ), .IN3(\mem[30][29] ), .IN2(\mem[29][29] ), .IN4(\mem[31][29] ), .S0(n1441), .S1(n1465), .Q(n1391) );
  MUX41X1 U1639 ( .IN1(\mem[24][29] ), .IN3(\mem[26][29] ), .IN2(\mem[25][29] ), .IN4(\mem[27][29] ), .S0(n1443), .S1(n1465), .Q(n1392) );
  MUX41X1 U1640 ( .IN1(\mem[20][29] ), .IN3(\mem[22][29] ), .IN2(\mem[21][29] ), .IN4(\mem[23][29] ), .S0(n1444), .S1(n1465), .Q(n1393) );
  MUX41X1 U1641 ( .IN1(\mem[16][29] ), .IN3(\mem[18][29] ), .IN2(\mem[17][29] ), .IN4(\mem[19][29] ), .S0(n1442), .S1(n1465), .Q(n1394) );
  MUX41X1 U1642 ( .IN1(n1394), .IN3(n1392), .IN2(n1393), .IN4(n1391), .S0(N13), 
        .S1(n1422), .Q(n1395) );
  MUX41X1 U1643 ( .IN1(\mem[12][29] ), .IN3(\mem[14][29] ), .IN2(\mem[13][29] ), .IN4(\mem[15][29] ), .S0(n1437), .S1(n1465), .Q(n1396) );
  MUX41X1 U1644 ( .IN1(\mem[8][29] ), .IN3(\mem[10][29] ), .IN2(\mem[9][29] ), 
        .IN4(\mem[11][29] ), .S0(n1440), .S1(n1465), .Q(n1397) );
  MUX41X1 U1645 ( .IN1(\mem[4][29] ), .IN3(\mem[6][29] ), .IN2(\mem[5][29] ), 
        .IN4(\mem[7][29] ), .S0(n1442), .S1(n1465), .Q(n1398) );
  MUX41X1 U1646 ( .IN1(\mem[0][29] ), .IN3(\mem[2][29] ), .IN2(\mem[1][29] ), 
        .IN4(\mem[3][29] ), .S0(n1441), .S1(n1465), .Q(n1399) );
  MUX41X1 U1647 ( .IN1(n1399), .IN3(n1397), .IN2(n1398), .IN4(n1396), .S0(N13), 
        .S1(n1422), .Q(n1400) );
  MUX21X1 U1648 ( .IN1(n1400), .IN2(n1395), .S(N14), .Q(rd_dataA[29]) );
  MUX41X1 U1649 ( .IN1(\mem[28][30] ), .IN3(\mem[30][30] ), .IN2(\mem[29][30] ), .IN4(\mem[31][30] ), .S0(N11), .S1(n1465), .Q(n1401) );
  MUX41X1 U1650 ( .IN1(\mem[24][30] ), .IN3(\mem[26][30] ), .IN2(\mem[25][30] ), .IN4(\mem[27][30] ), .S0(n1444), .S1(n1465), .Q(n1402) );
  MUX41X1 U1651 ( .IN1(\mem[20][30] ), .IN3(\mem[22][30] ), .IN2(\mem[21][30] ), .IN4(\mem[23][30] ), .S0(n1440), .S1(n1465), .Q(n1403) );
  MUX41X1 U1652 ( .IN1(\mem[16][30] ), .IN3(\mem[18][30] ), .IN2(\mem[17][30] ), .IN4(\mem[19][30] ), .S0(n1443), .S1(n1465), .Q(n1404) );
  MUX41X1 U1653 ( .IN1(n1404), .IN3(n1402), .IN2(n1403), .IN4(n1401), .S0(N13), 
        .S1(n1422), .Q(n1405) );
  MUX41X1 U1654 ( .IN1(\mem[12][30] ), .IN3(\mem[14][30] ), .IN2(\mem[13][30] ), .IN4(\mem[15][30] ), .S0(N11), .S1(n1460), .Q(n1406) );
  MUX41X1 U1655 ( .IN1(\mem[8][30] ), .IN3(\mem[10][30] ), .IN2(\mem[9][30] ), 
        .IN4(\mem[11][30] ), .S0(N11), .S1(n1457), .Q(n1407) );
  MUX41X1 U1656 ( .IN1(\mem[4][30] ), .IN3(\mem[6][30] ), .IN2(\mem[5][30] ), 
        .IN4(\mem[7][30] ), .S0(n1442), .S1(N10), .Q(n1408) );
  MUX41X1 U1657 ( .IN1(\mem[0][30] ), .IN3(\mem[2][30] ), .IN2(\mem[1][30] ), 
        .IN4(\mem[3][30] ), .S0(n1440), .S1(n1465), .Q(n1409) );
  MUX41X1 U1658 ( .IN1(n1409), .IN3(n1407), .IN2(n1408), .IN4(n1406), .S0(N13), 
        .S1(N12), .Q(n1410) );
  MUX21X1 U1659 ( .IN1(n1410), .IN2(n1405), .S(N14), .Q(rd_dataA[30]) );
  MUX41X1 U1660 ( .IN1(\mem[28][31] ), .IN3(\mem[30][31] ), .IN2(\mem[29][31] ), .IN4(\mem[31][31] ), .S0(N11), .S1(n1459), .Q(n1411) );
  MUX41X1 U1661 ( .IN1(\mem[24][31] ), .IN3(\mem[26][31] ), .IN2(\mem[25][31] ), .IN4(\mem[27][31] ), .S0(n1444), .S1(N10), .Q(n1412) );
  MUX41X1 U1662 ( .IN1(\mem[20][31] ), .IN3(\mem[22][31] ), .IN2(\mem[21][31] ), .IN4(\mem[23][31] ), .S0(n1439), .S1(n1464), .Q(n1413) );
  MUX41X1 U1663 ( .IN1(\mem[16][31] ), .IN3(\mem[18][31] ), .IN2(\mem[17][31] ), .IN4(\mem[19][31] ), .S0(n1437), .S1(n1462), .Q(n1414) );
  MUX41X1 U1664 ( .IN1(n1414), .IN3(n1412), .IN2(n1413), .IN4(n1411), .S0(N13), 
        .S1(n1423), .Q(n1415) );
  MUX41X1 U1665 ( .IN1(\mem[12][31] ), .IN3(\mem[14][31] ), .IN2(\mem[13][31] ), .IN4(\mem[15][31] ), .S0(N11), .S1(n1461), .Q(n1416) );
  MUX41X1 U1666 ( .IN1(\mem[8][31] ), .IN3(\mem[10][31] ), .IN2(\mem[9][31] ), 
        .IN4(\mem[11][31] ), .S0(N11), .S1(n1458), .Q(n1417) );
  MUX41X1 U1667 ( .IN1(\mem[4][31] ), .IN3(\mem[6][31] ), .IN2(\mem[5][31] ), 
        .IN4(\mem[7][31] ), .S0(n1443), .S1(N10), .Q(n1418) );
  MUX41X1 U1668 ( .IN1(\mem[0][31] ), .IN3(\mem[2][31] ), .IN2(\mem[1][31] ), 
        .IN4(\mem[3][31] ), .S0(n1441), .S1(N10), .Q(n1419) );
  MUX41X1 U1669 ( .IN1(n1419), .IN3(n1417), .IN2(n1418), .IN4(n1416), .S0(N13), 
        .S1(N12), .Q(n1420) );
  MUX21X1 U1670 ( .IN1(n1420), .IN2(n1415), .S(N14), .Q(rd_dataA[31]) );
  MUX41X1 U1671 ( .IN1(\mem[28][0] ), .IN3(\mem[30][0] ), .IN2(\mem[29][0] ), 
        .IN4(\mem[31][0] ), .S0(n1810), .S1(n1822), .Q(n1466) );
  MUX41X1 U1672 ( .IN1(\mem[24][0] ), .IN3(\mem[26][0] ), .IN2(\mem[25][0] ), 
        .IN4(\mem[27][0] ), .S0(n1809), .S1(n1821), .Q(n1467) );
  MUX41X1 U1673 ( .IN1(\mem[20][0] ), .IN3(\mem[22][0] ), .IN2(\mem[21][0] ), 
        .IN4(\mem[23][0] ), .S0(n1807), .S1(n1819), .Q(n1468) );
  MUX41X1 U1674 ( .IN1(\mem[16][0] ), .IN3(\mem[18][0] ), .IN2(\mem[17][0] ), 
        .IN4(\mem[19][0] ), .S0(n1811), .S1(n1818), .Q(n1469) );
  MUX41X1 U1675 ( .IN1(n1469), .IN3(n1467), .IN2(n1468), .IN4(n1466), .S0(N18), 
        .S1(n1790), .Q(n1470) );
  MUX41X1 U1676 ( .IN1(\mem[12][0] ), .IN3(\mem[14][0] ), .IN2(\mem[13][0] ), 
        .IN4(\mem[15][0] ), .S0(n1793), .S1(n1814), .Q(n1471) );
  MUX41X1 U1677 ( .IN1(\mem[8][0] ), .IN3(\mem[10][0] ), .IN2(\mem[9][0] ), 
        .IN4(\mem[11][0] ), .S0(n1793), .S1(n1814), .Q(n1472) );
  MUX41X1 U1678 ( .IN1(\mem[4][0] ), .IN3(\mem[6][0] ), .IN2(\mem[5][0] ), 
        .IN4(\mem[7][0] ), .S0(n1793), .S1(n1814), .Q(n1473) );
  MUX41X1 U1679 ( .IN1(\mem[0][0] ), .IN3(\mem[2][0] ), .IN2(\mem[1][0] ), 
        .IN4(\mem[3][0] ), .S0(n1793), .S1(n1814), .Q(n1474) );
  MUX41X1 U1680 ( .IN1(n1474), .IN3(n1472), .IN2(n1473), .IN4(n1471), .S0(N18), 
        .S1(n1790), .Q(n1475) );
  MUX21X1 U1681 ( .IN1(n1475), .IN2(n1470), .S(N19), .Q(rd_dataB[0]) );
  MUX41X1 U1682 ( .IN1(\mem[28][1] ), .IN3(\mem[30][1] ), .IN2(\mem[29][1] ), 
        .IN4(\mem[31][1] ), .S0(n1793), .S1(n1814), .Q(n1476) );
  MUX41X1 U1683 ( .IN1(\mem[24][1] ), .IN3(\mem[26][1] ), .IN2(\mem[25][1] ), 
        .IN4(\mem[27][1] ), .S0(n1793), .S1(n1814), .Q(n1477) );
  MUX41X1 U1684 ( .IN1(\mem[20][1] ), .IN3(\mem[22][1] ), .IN2(\mem[21][1] ), 
        .IN4(\mem[23][1] ), .S0(n1793), .S1(n1814), .Q(n1478) );
  MUX41X1 U1685 ( .IN1(\mem[16][1] ), .IN3(\mem[18][1] ), .IN2(\mem[17][1] ), 
        .IN4(\mem[19][1] ), .S0(n1793), .S1(n1814), .Q(n1479) );
  MUX41X1 U1686 ( .IN1(n1479), .IN3(n1477), .IN2(n1478), .IN4(n1476), .S0(N18), 
        .S1(n1790), .Q(n1480) );
  MUX41X1 U1687 ( .IN1(\mem[12][1] ), .IN3(\mem[14][1] ), .IN2(\mem[13][1] ), 
        .IN4(\mem[15][1] ), .S0(n1793), .S1(n1814), .Q(n1481) );
  MUX41X1 U1688 ( .IN1(\mem[8][1] ), .IN3(\mem[10][1] ), .IN2(\mem[9][1] ), 
        .IN4(\mem[11][1] ), .S0(n1793), .S1(n1814), .Q(n1482) );
  MUX41X1 U1689 ( .IN1(\mem[4][1] ), .IN3(\mem[6][1] ), .IN2(\mem[5][1] ), 
        .IN4(\mem[7][1] ), .S0(n1793), .S1(n1814), .Q(n1483) );
  MUX41X1 U1690 ( .IN1(\mem[0][1] ), .IN3(\mem[2][1] ), .IN2(\mem[1][1] ), 
        .IN4(\mem[3][1] ), .S0(n1793), .S1(n1814), .Q(n1484) );
  MUX41X1 U1691 ( .IN1(n1484), .IN3(n1482), .IN2(n1483), .IN4(n1481), .S0(N18), 
        .S1(n1790), .Q(n1485) );
  MUX21X1 U1692 ( .IN1(n1485), .IN2(n1480), .S(N19), .Q(rd_dataB[1]) );
  MUX41X1 U1693 ( .IN1(\mem[28][2] ), .IN3(\mem[30][2] ), .IN2(\mem[29][2] ), 
        .IN4(\mem[31][2] ), .S0(n1794), .S1(n1815), .Q(n1486) );
  MUX41X1 U1694 ( .IN1(\mem[24][2] ), .IN3(\mem[26][2] ), .IN2(\mem[25][2] ), 
        .IN4(\mem[27][2] ), .S0(n1794), .S1(n1815), .Q(n1487) );
  MUX41X1 U1695 ( .IN1(\mem[20][2] ), .IN3(\mem[22][2] ), .IN2(\mem[21][2] ), 
        .IN4(\mem[23][2] ), .S0(n1794), .S1(n1815), .Q(n1488) );
  MUX41X1 U1696 ( .IN1(\mem[16][2] ), .IN3(\mem[18][2] ), .IN2(\mem[17][2] ), 
        .IN4(\mem[19][2] ), .S0(n1794), .S1(n1815), .Q(n1489) );
  MUX41X1 U1697 ( .IN1(n1489), .IN3(n1487), .IN2(n1488), .IN4(n1486), .S0(N18), 
        .S1(n1790), .Q(n1490) );
  MUX41X1 U1698 ( .IN1(\mem[12][2] ), .IN3(\mem[14][2] ), .IN2(\mem[13][2] ), 
        .IN4(\mem[15][2] ), .S0(n1794), .S1(n1815), .Q(n1491) );
  MUX41X1 U1699 ( .IN1(\mem[8][2] ), .IN3(\mem[10][2] ), .IN2(\mem[9][2] ), 
        .IN4(\mem[11][2] ), .S0(n1794), .S1(n1815), .Q(n1492) );
  MUX41X1 U1700 ( .IN1(\mem[4][2] ), .IN3(\mem[6][2] ), .IN2(\mem[5][2] ), 
        .IN4(\mem[7][2] ), .S0(n1794), .S1(n1815), .Q(n1493) );
  MUX41X1 U1701 ( .IN1(\mem[0][2] ), .IN3(\mem[2][2] ), .IN2(\mem[1][2] ), 
        .IN4(\mem[3][2] ), .S0(n1794), .S1(n1815), .Q(n1494) );
  MUX41X1 U1702 ( .IN1(n1494), .IN3(n1492), .IN2(n1493), .IN4(n1491), .S0(N18), 
        .S1(n1790), .Q(n1495) );
  MUX21X1 U1703 ( .IN1(n1495), .IN2(n1490), .S(N19), .Q(rd_dataB[2]) );
  MUX41X1 U1704 ( .IN1(\mem[28][3] ), .IN3(\mem[30][3] ), .IN2(\mem[29][3] ), 
        .IN4(\mem[31][3] ), .S0(n1794), .S1(n1815), .Q(n1496) );
  MUX41X1 U1705 ( .IN1(\mem[24][3] ), .IN3(\mem[26][3] ), .IN2(\mem[25][3] ), 
        .IN4(\mem[27][3] ), .S0(n1794), .S1(n1815), .Q(n1497) );
  MUX41X1 U1706 ( .IN1(\mem[20][3] ), .IN3(\mem[22][3] ), .IN2(\mem[21][3] ), 
        .IN4(\mem[23][3] ), .S0(n1794), .S1(n1815), .Q(n1498) );
  MUX41X1 U1707 ( .IN1(\mem[16][3] ), .IN3(\mem[18][3] ), .IN2(\mem[17][3] ), 
        .IN4(\mem[19][3] ), .S0(n1794), .S1(n1815), .Q(n1499) );
  MUX41X1 U1708 ( .IN1(n1499), .IN3(n1497), .IN2(n1498), .IN4(n1496), .S0(N18), 
        .S1(n1790), .Q(n1500) );
  MUX41X1 U1709 ( .IN1(\mem[12][3] ), .IN3(\mem[14][3] ), .IN2(\mem[13][3] ), 
        .IN4(\mem[15][3] ), .S0(n1795), .S1(n1816), .Q(n1501) );
  MUX41X1 U1710 ( .IN1(\mem[8][3] ), .IN3(\mem[10][3] ), .IN2(\mem[9][3] ), 
        .IN4(\mem[11][3] ), .S0(n1795), .S1(n1816), .Q(n1502) );
  MUX41X1 U1711 ( .IN1(\mem[4][3] ), .IN3(\mem[6][3] ), .IN2(\mem[5][3] ), 
        .IN4(\mem[7][3] ), .S0(n1795), .S1(n1816), .Q(n1503) );
  MUX41X1 U1712 ( .IN1(\mem[0][3] ), .IN3(\mem[2][3] ), .IN2(\mem[1][3] ), 
        .IN4(\mem[3][3] ), .S0(n1795), .S1(n1816), .Q(n1504) );
  MUX41X1 U1713 ( .IN1(n1504), .IN3(n1502), .IN2(n1503), .IN4(n1501), .S0(N18), 
        .S1(n1790), .Q(n1505) );
  MUX21X1 U1714 ( .IN1(n1505), .IN2(n1500), .S(N19), .Q(rd_dataB[3]) );
  MUX41X1 U1715 ( .IN1(\mem[28][4] ), .IN3(\mem[30][4] ), .IN2(\mem[29][4] ), 
        .IN4(\mem[31][4] ), .S0(n1795), .S1(n1816), .Q(n1506) );
  MUX41X1 U1716 ( .IN1(\mem[24][4] ), .IN3(\mem[26][4] ), .IN2(\mem[25][4] ), 
        .IN4(\mem[27][4] ), .S0(n1795), .S1(n1816), .Q(n1507) );
  MUX41X1 U1717 ( .IN1(\mem[20][4] ), .IN3(\mem[22][4] ), .IN2(\mem[21][4] ), 
        .IN4(\mem[23][4] ), .S0(n1795), .S1(n1816), .Q(n1508) );
  MUX41X1 U1718 ( .IN1(\mem[16][4] ), .IN3(\mem[18][4] ), .IN2(\mem[17][4] ), 
        .IN4(\mem[19][4] ), .S0(n1795), .S1(n1816), .Q(n1509) );
  MUX41X1 U1719 ( .IN1(n1509), .IN3(n1507), .IN2(n1508), .IN4(n1506), .S0(N18), 
        .S1(n1790), .Q(n1510) );
  MUX41X1 U1720 ( .IN1(\mem[12][4] ), .IN3(\mem[14][4] ), .IN2(\mem[13][4] ), 
        .IN4(\mem[15][4] ), .S0(n1795), .S1(n1816), .Q(n1511) );
  MUX41X1 U1721 ( .IN1(\mem[8][4] ), .IN3(\mem[10][4] ), .IN2(\mem[9][4] ), 
        .IN4(\mem[11][4] ), .S0(n1795), .S1(n1816), .Q(n1512) );
  MUX41X1 U1722 ( .IN1(\mem[4][4] ), .IN3(\mem[6][4] ), .IN2(\mem[5][4] ), 
        .IN4(\mem[7][4] ), .S0(n1795), .S1(n1816), .Q(n1513) );
  MUX41X1 U1723 ( .IN1(\mem[0][4] ), .IN3(\mem[2][4] ), .IN2(\mem[1][4] ), 
        .IN4(\mem[3][4] ), .S0(n1795), .S1(n1816), .Q(n1514) );
  MUX41X1 U1724 ( .IN1(n1514), .IN3(n1512), .IN2(n1513), .IN4(n1511), .S0(N18), 
        .S1(n1790), .Q(n1515) );
  MUX21X1 U1725 ( .IN1(n1515), .IN2(n1510), .S(N19), .Q(rd_dataB[4]) );
  MUX41X1 U1726 ( .IN1(\mem[28][5] ), .IN3(\mem[30][5] ), .IN2(\mem[29][5] ), 
        .IN4(\mem[31][5] ), .S0(n1796), .S1(n1817), .Q(n1516) );
  MUX41X1 U1727 ( .IN1(\mem[24][5] ), .IN3(\mem[26][5] ), .IN2(\mem[25][5] ), 
        .IN4(\mem[27][5] ), .S0(n1796), .S1(n1817), .Q(n1517) );
  MUX41X1 U1728 ( .IN1(\mem[20][5] ), .IN3(\mem[22][5] ), .IN2(\mem[21][5] ), 
        .IN4(\mem[23][5] ), .S0(n1796), .S1(n1817), .Q(n1518) );
  MUX41X1 U1729 ( .IN1(\mem[16][5] ), .IN3(\mem[18][5] ), .IN2(\mem[17][5] ), 
        .IN4(\mem[19][5] ), .S0(n1796), .S1(n1817), .Q(n1519) );
  MUX41X1 U1730 ( .IN1(n1519), .IN3(n1517), .IN2(n1518), .IN4(n1516), .S0(N18), 
        .S1(n1790), .Q(n1520) );
  MUX41X1 U1731 ( .IN1(\mem[12][5] ), .IN3(\mem[14][5] ), .IN2(\mem[13][5] ), 
        .IN4(\mem[15][5] ), .S0(n1796), .S1(n1817), .Q(n1521) );
  MUX41X1 U1732 ( .IN1(\mem[8][5] ), .IN3(\mem[10][5] ), .IN2(\mem[9][5] ), 
        .IN4(\mem[11][5] ), .S0(n1796), .S1(n1817), .Q(n1522) );
  MUX41X1 U1733 ( .IN1(\mem[4][5] ), .IN3(\mem[6][5] ), .IN2(\mem[5][5] ), 
        .IN4(\mem[7][5] ), .S0(n1796), .S1(n1817), .Q(n1523) );
  MUX41X1 U1734 ( .IN1(\mem[0][5] ), .IN3(\mem[2][5] ), .IN2(\mem[1][5] ), 
        .IN4(\mem[3][5] ), .S0(n1796), .S1(n1817), .Q(n1524) );
  MUX41X1 U1735 ( .IN1(n1524), .IN3(n1522), .IN2(n1523), .IN4(n1521), .S0(N18), 
        .S1(n1790), .Q(n1525) );
  MUX21X1 U1736 ( .IN1(n1525), .IN2(n1520), .S(N19), .Q(rd_dataB[5]) );
  MUX41X1 U1737 ( .IN1(\mem[28][6] ), .IN3(\mem[30][6] ), .IN2(\mem[29][6] ), 
        .IN4(\mem[31][6] ), .S0(n1796), .S1(n1817), .Q(n1526) );
  MUX41X1 U1738 ( .IN1(\mem[24][6] ), .IN3(\mem[26][6] ), .IN2(\mem[25][6] ), 
        .IN4(\mem[27][6] ), .S0(n1796), .S1(n1817), .Q(n1527) );
  MUX41X1 U1739 ( .IN1(\mem[20][6] ), .IN3(\mem[22][6] ), .IN2(\mem[21][6] ), 
        .IN4(\mem[23][6] ), .S0(n1796), .S1(n1817), .Q(n1528) );
  MUX41X1 U1740 ( .IN1(\mem[16][6] ), .IN3(\mem[18][6] ), .IN2(\mem[17][6] ), 
        .IN4(\mem[19][6] ), .S0(n1796), .S1(n1817), .Q(n1529) );
  MUX41X1 U1741 ( .IN1(n1529), .IN3(n1527), .IN2(n1528), .IN4(n1526), .S0(N18), 
        .S1(n1789), .Q(n1530) );
  MUX41X1 U1742 ( .IN1(\mem[12][6] ), .IN3(\mem[14][6] ), .IN2(\mem[13][6] ), 
        .IN4(\mem[15][6] ), .S0(n1797), .S1(n1818), .Q(n1531) );
  MUX41X1 U1743 ( .IN1(\mem[8][6] ), .IN3(\mem[10][6] ), .IN2(\mem[9][6] ), 
        .IN4(\mem[11][6] ), .S0(n1797), .S1(n1818), .Q(n1532) );
  MUX41X1 U1744 ( .IN1(\mem[4][6] ), .IN3(\mem[6][6] ), .IN2(\mem[5][6] ), 
        .IN4(\mem[7][6] ), .S0(n1797), .S1(n1818), .Q(n1533) );
  MUX41X1 U1745 ( .IN1(\mem[0][6] ), .IN3(\mem[2][6] ), .IN2(\mem[1][6] ), 
        .IN4(\mem[3][6] ), .S0(n1797), .S1(n1818), .Q(n1534) );
  MUX41X1 U1746 ( .IN1(n1534), .IN3(n1532), .IN2(n1533), .IN4(n1531), .S0(N18), 
        .S1(n1789), .Q(n1535) );
  MUX21X1 U1747 ( .IN1(n1535), .IN2(n1530), .S(N19), .Q(rd_dataB[6]) );
  MUX41X1 U1748 ( .IN1(\mem[28][7] ), .IN3(\mem[30][7] ), .IN2(\mem[29][7] ), 
        .IN4(\mem[31][7] ), .S0(n1797), .S1(n1818), .Q(n1536) );
  MUX41X1 U1749 ( .IN1(\mem[24][7] ), .IN3(\mem[26][7] ), .IN2(\mem[25][7] ), 
        .IN4(\mem[27][7] ), .S0(n1797), .S1(n1818), .Q(n1537) );
  MUX41X1 U1750 ( .IN1(\mem[20][7] ), .IN3(\mem[22][7] ), .IN2(\mem[21][7] ), 
        .IN4(\mem[23][7] ), .S0(n1797), .S1(n1818), .Q(n1538) );
  MUX41X1 U1751 ( .IN1(\mem[16][7] ), .IN3(\mem[18][7] ), .IN2(\mem[17][7] ), 
        .IN4(\mem[19][7] ), .S0(n1797), .S1(n1818), .Q(n1539) );
  MUX41X1 U1752 ( .IN1(n1539), .IN3(n1537), .IN2(n1538), .IN4(n1536), .S0(N18), 
        .S1(n1789), .Q(n1540) );
  MUX41X1 U1753 ( .IN1(\mem[12][7] ), .IN3(\mem[14][7] ), .IN2(\mem[13][7] ), 
        .IN4(\mem[15][7] ), .S0(n1797), .S1(n1818), .Q(n1541) );
  MUX41X1 U1754 ( .IN1(\mem[8][7] ), .IN3(\mem[10][7] ), .IN2(\mem[9][7] ), 
        .IN4(\mem[11][7] ), .S0(n1797), .S1(n1818), .Q(n1542) );
  MUX41X1 U1755 ( .IN1(\mem[4][7] ), .IN3(\mem[6][7] ), .IN2(\mem[5][7] ), 
        .IN4(\mem[7][7] ), .S0(n1797), .S1(n1818), .Q(n1543) );
  MUX41X1 U1756 ( .IN1(\mem[0][7] ), .IN3(\mem[2][7] ), .IN2(\mem[1][7] ), 
        .IN4(\mem[3][7] ), .S0(n1797), .S1(n1818), .Q(n1544) );
  MUX41X1 U1757 ( .IN1(n1544), .IN3(n1542), .IN2(n1543), .IN4(n1541), .S0(N18), 
        .S1(n1789), .Q(n1545) );
  MUX21X1 U1758 ( .IN1(n1545), .IN2(n1540), .S(N19), .Q(rd_dataB[7]) );
  MUX41X1 U1759 ( .IN1(\mem[28][8] ), .IN3(\mem[30][8] ), .IN2(\mem[29][8] ), 
        .IN4(\mem[31][8] ), .S0(n1798), .S1(n1819), .Q(n1546) );
  MUX41X1 U1760 ( .IN1(\mem[24][8] ), .IN3(\mem[26][8] ), .IN2(\mem[25][8] ), 
        .IN4(\mem[27][8] ), .S0(n1798), .S1(n1819), .Q(n1547) );
  MUX41X1 U1761 ( .IN1(\mem[20][8] ), .IN3(\mem[22][8] ), .IN2(\mem[21][8] ), 
        .IN4(\mem[23][8] ), .S0(n1798), .S1(n1819), .Q(n1548) );
  MUX41X1 U1762 ( .IN1(\mem[16][8] ), .IN3(\mem[18][8] ), .IN2(\mem[17][8] ), 
        .IN4(\mem[19][8] ), .S0(n1798), .S1(n1819), .Q(n1549) );
  MUX41X1 U1763 ( .IN1(n1549), .IN3(n1547), .IN2(n1548), .IN4(n1546), .S0(N18), 
        .S1(n1789), .Q(n1550) );
  MUX41X1 U1764 ( .IN1(\mem[12][8] ), .IN3(\mem[14][8] ), .IN2(\mem[13][8] ), 
        .IN4(\mem[15][8] ), .S0(n1798), .S1(n1819), .Q(n1551) );
  MUX41X1 U1765 ( .IN1(\mem[8][8] ), .IN3(\mem[10][8] ), .IN2(\mem[9][8] ), 
        .IN4(\mem[11][8] ), .S0(n1798), .S1(n1819), .Q(n1552) );
  MUX41X1 U1766 ( .IN1(\mem[4][8] ), .IN3(\mem[6][8] ), .IN2(\mem[5][8] ), 
        .IN4(\mem[7][8] ), .S0(n1798), .S1(n1819), .Q(n1553) );
  MUX41X1 U1767 ( .IN1(\mem[0][8] ), .IN3(\mem[2][8] ), .IN2(\mem[1][8] ), 
        .IN4(\mem[3][8] ), .S0(n1798), .S1(n1819), .Q(n1554) );
  MUX41X1 U1768 ( .IN1(n1554), .IN3(n1552), .IN2(n1553), .IN4(n1551), .S0(N18), 
        .S1(n1789), .Q(n1555) );
  MUX21X1 U1769 ( .IN1(n1555), .IN2(n1550), .S(N19), .Q(rd_dataB[8]) );
  MUX41X1 U1770 ( .IN1(\mem[28][9] ), .IN3(\mem[30][9] ), .IN2(\mem[29][9] ), 
        .IN4(\mem[31][9] ), .S0(n1798), .S1(n1819), .Q(n1556) );
  MUX41X1 U1771 ( .IN1(\mem[24][9] ), .IN3(\mem[26][9] ), .IN2(\mem[25][9] ), 
        .IN4(\mem[27][9] ), .S0(n1798), .S1(n1819), .Q(n1557) );
  MUX41X1 U1772 ( .IN1(\mem[20][9] ), .IN3(\mem[22][9] ), .IN2(\mem[21][9] ), 
        .IN4(\mem[23][9] ), .S0(n1798), .S1(n1819), .Q(n1558) );
  MUX41X1 U1773 ( .IN1(\mem[16][9] ), .IN3(\mem[18][9] ), .IN2(\mem[17][9] ), 
        .IN4(\mem[19][9] ), .S0(n1798), .S1(n1819), .Q(n1559) );
  MUX41X1 U1774 ( .IN1(n1559), .IN3(n1557), .IN2(n1558), .IN4(n1556), .S0(N18), 
        .S1(n1789), .Q(n1560) );
  MUX41X1 U1775 ( .IN1(\mem[12][9] ), .IN3(\mem[14][9] ), .IN2(\mem[13][9] ), 
        .IN4(\mem[15][9] ), .S0(n1799), .S1(n1820), .Q(n1561) );
  MUX41X1 U1776 ( .IN1(\mem[8][9] ), .IN3(\mem[10][9] ), .IN2(\mem[9][9] ), 
        .IN4(\mem[11][9] ), .S0(n1799), .S1(n1820), .Q(n1562) );
  MUX41X1 U1777 ( .IN1(\mem[4][9] ), .IN3(\mem[6][9] ), .IN2(\mem[5][9] ), 
        .IN4(\mem[7][9] ), .S0(n1799), .S1(n1820), .Q(n1563) );
  MUX41X1 U1778 ( .IN1(\mem[0][9] ), .IN3(\mem[2][9] ), .IN2(\mem[1][9] ), 
        .IN4(\mem[3][9] ), .S0(n1799), .S1(n1820), .Q(n1564) );
  MUX41X1 U1779 ( .IN1(n1564), .IN3(n1562), .IN2(n1563), .IN4(n1561), .S0(N18), 
        .S1(n1789), .Q(n1565) );
  MUX21X1 U1780 ( .IN1(n1565), .IN2(n1560), .S(N19), .Q(rd_dataB[9]) );
  MUX41X1 U1781 ( .IN1(\mem[28][10] ), .IN3(\mem[30][10] ), .IN2(\mem[29][10] ), .IN4(\mem[31][10] ), .S0(n1799), .S1(n1820), .Q(n1566) );
  MUX41X1 U1782 ( .IN1(\mem[24][10] ), .IN3(\mem[26][10] ), .IN2(\mem[25][10] ), .IN4(\mem[27][10] ), .S0(n1799), .S1(n1820), .Q(n1567) );
  MUX41X1 U1783 ( .IN1(\mem[20][10] ), .IN3(\mem[22][10] ), .IN2(\mem[21][10] ), .IN4(\mem[23][10] ), .S0(n1799), .S1(n1820), .Q(n1568) );
  MUX41X1 U1784 ( .IN1(\mem[16][10] ), .IN3(\mem[18][10] ), .IN2(\mem[17][10] ), .IN4(\mem[19][10] ), .S0(n1799), .S1(n1820), .Q(n1569) );
  MUX41X1 U1785 ( .IN1(n1569), .IN3(n1567), .IN2(n1568), .IN4(n1566), .S0(N18), 
        .S1(n1789), .Q(n1570) );
  MUX41X1 U1786 ( .IN1(\mem[12][10] ), .IN3(\mem[14][10] ), .IN2(\mem[13][10] ), .IN4(\mem[15][10] ), .S0(n1799), .S1(n1820), .Q(n1571) );
  MUX41X1 U1787 ( .IN1(\mem[8][10] ), .IN3(\mem[10][10] ), .IN2(\mem[9][10] ), 
        .IN4(\mem[11][10] ), .S0(n1799), .S1(n1820), .Q(n1572) );
  MUX41X1 U1788 ( .IN1(\mem[4][10] ), .IN3(\mem[6][10] ), .IN2(\mem[5][10] ), 
        .IN4(\mem[7][10] ), .S0(n1799), .S1(n1820), .Q(n1573) );
  MUX41X1 U1789 ( .IN1(\mem[0][10] ), .IN3(\mem[2][10] ), .IN2(\mem[1][10] ), 
        .IN4(\mem[3][10] ), .S0(n1799), .S1(n1820), .Q(n1574) );
  MUX41X1 U1790 ( .IN1(n1574), .IN3(n1572), .IN2(n1573), .IN4(n1571), .S0(N18), 
        .S1(n1789), .Q(n1575) );
  MUX21X1 U1791 ( .IN1(n1575), .IN2(n1570), .S(N19), .Q(rd_dataB[10]) );
  MUX41X1 U1792 ( .IN1(\mem[28][11] ), .IN3(\mem[30][11] ), .IN2(\mem[29][11] ), .IN4(\mem[31][11] ), .S0(n1800), .S1(n1821), .Q(n1576) );
  MUX41X1 U1793 ( .IN1(\mem[24][11] ), .IN3(\mem[26][11] ), .IN2(\mem[25][11] ), .IN4(\mem[27][11] ), .S0(n1800), .S1(n1821), .Q(n1577) );
  MUX41X1 U1794 ( .IN1(\mem[20][11] ), .IN3(\mem[22][11] ), .IN2(\mem[21][11] ), .IN4(\mem[23][11] ), .S0(n1800), .S1(n1821), .Q(n1578) );
  MUX41X1 U1795 ( .IN1(\mem[16][11] ), .IN3(\mem[18][11] ), .IN2(\mem[17][11] ), .IN4(\mem[19][11] ), .S0(n1800), .S1(n1821), .Q(n1579) );
  MUX41X1 U1796 ( .IN1(n1579), .IN3(n1577), .IN2(n1578), .IN4(n1576), .S0(N18), 
        .S1(n1789), .Q(n1580) );
  MUX41X1 U1797 ( .IN1(\mem[12][11] ), .IN3(\mem[14][11] ), .IN2(\mem[13][11] ), .IN4(\mem[15][11] ), .S0(n1800), .S1(n1821), .Q(n1581) );
  MUX41X1 U1798 ( .IN1(\mem[8][11] ), .IN3(\mem[10][11] ), .IN2(\mem[9][11] ), 
        .IN4(\mem[11][11] ), .S0(n1800), .S1(n1821), .Q(n1582) );
  MUX41X1 U1799 ( .IN1(\mem[4][11] ), .IN3(\mem[6][11] ), .IN2(\mem[5][11] ), 
        .IN4(\mem[7][11] ), .S0(n1800), .S1(n1821), .Q(n1583) );
  MUX41X1 U1800 ( .IN1(\mem[0][11] ), .IN3(\mem[2][11] ), .IN2(\mem[1][11] ), 
        .IN4(\mem[3][11] ), .S0(n1800), .S1(n1821), .Q(n1584) );
  MUX41X1 U1801 ( .IN1(n1584), .IN3(n1582), .IN2(n1583), .IN4(n1581), .S0(N18), 
        .S1(n1789), .Q(n1585) );
  MUX21X1 U1802 ( .IN1(n1585), .IN2(n1580), .S(N19), .Q(rd_dataB[11]) );
  MUX41X1 U1803 ( .IN1(\mem[28][12] ), .IN3(\mem[30][12] ), .IN2(\mem[29][12] ), .IN4(\mem[31][12] ), .S0(n1800), .S1(n1821), .Q(n1586) );
  MUX41X1 U1804 ( .IN1(\mem[24][12] ), .IN3(\mem[26][12] ), .IN2(\mem[25][12] ), .IN4(\mem[27][12] ), .S0(n1800), .S1(n1821), .Q(n1587) );
  MUX41X1 U1805 ( .IN1(\mem[20][12] ), .IN3(\mem[22][12] ), .IN2(\mem[21][12] ), .IN4(\mem[23][12] ), .S0(n1800), .S1(n1821), .Q(n1588) );
  MUX41X1 U1806 ( .IN1(\mem[16][12] ), .IN3(\mem[18][12] ), .IN2(\mem[17][12] ), .IN4(\mem[19][12] ), .S0(n1800), .S1(n1821), .Q(n1589) );
  MUX41X1 U1807 ( .IN1(n1589), .IN3(n1587), .IN2(n1588), .IN4(n1586), .S0(N18), 
        .S1(n1788), .Q(n1590) );
  MUX41X1 U1808 ( .IN1(\mem[12][12] ), .IN3(\mem[14][12] ), .IN2(\mem[13][12] ), .IN4(\mem[15][12] ), .S0(n1801), .S1(n1822), .Q(n1591) );
  MUX41X1 U1809 ( .IN1(\mem[8][12] ), .IN3(\mem[10][12] ), .IN2(\mem[9][12] ), 
        .IN4(\mem[11][12] ), .S0(n1801), .S1(n1822), .Q(n1592) );
  MUX41X1 U1810 ( .IN1(\mem[4][12] ), .IN3(\mem[6][12] ), .IN2(\mem[5][12] ), 
        .IN4(\mem[7][12] ), .S0(n1801), .S1(n1822), .Q(n1593) );
  MUX41X1 U1811 ( .IN1(\mem[0][12] ), .IN3(\mem[2][12] ), .IN2(\mem[1][12] ), 
        .IN4(\mem[3][12] ), .S0(n1801), .S1(n1822), .Q(n1594) );
  MUX41X1 U1812 ( .IN1(n1594), .IN3(n1592), .IN2(n1593), .IN4(n1591), .S0(N18), 
        .S1(n1788), .Q(n1595) );
  MUX21X1 U1813 ( .IN1(n1595), .IN2(n1590), .S(N19), .Q(rd_dataB[12]) );
  MUX41X1 U1814 ( .IN1(\mem[28][13] ), .IN3(\mem[30][13] ), .IN2(\mem[29][13] ), .IN4(\mem[31][13] ), .S0(n1801), .S1(n1822), .Q(n1596) );
  MUX41X1 U1815 ( .IN1(\mem[24][13] ), .IN3(\mem[26][13] ), .IN2(\mem[25][13] ), .IN4(\mem[27][13] ), .S0(n1801), .S1(n1822), .Q(n1597) );
  MUX41X1 U1816 ( .IN1(\mem[20][13] ), .IN3(\mem[22][13] ), .IN2(\mem[21][13] ), .IN4(\mem[23][13] ), .S0(n1801), .S1(n1822), .Q(n1598) );
  MUX41X1 U1817 ( .IN1(\mem[16][13] ), .IN3(\mem[18][13] ), .IN2(\mem[17][13] ), .IN4(\mem[19][13] ), .S0(n1801), .S1(n1822), .Q(n1599) );
  MUX41X1 U1818 ( .IN1(n1599), .IN3(n1597), .IN2(n1598), .IN4(n1596), .S0(N18), 
        .S1(n1788), .Q(n1600) );
  MUX41X1 U1819 ( .IN1(\mem[12][13] ), .IN3(\mem[14][13] ), .IN2(\mem[13][13] ), .IN4(\mem[15][13] ), .S0(n1801), .S1(n1822), .Q(n1601) );
  MUX41X1 U1820 ( .IN1(\mem[8][13] ), .IN3(\mem[10][13] ), .IN2(\mem[9][13] ), 
        .IN4(\mem[11][13] ), .S0(n1801), .S1(n1822), .Q(n1602) );
  MUX41X1 U1821 ( .IN1(\mem[4][13] ), .IN3(\mem[6][13] ), .IN2(\mem[5][13] ), 
        .IN4(\mem[7][13] ), .S0(n1801), .S1(n1822), .Q(n1603) );
  MUX41X1 U1822 ( .IN1(\mem[0][13] ), .IN3(\mem[2][13] ), .IN2(\mem[1][13] ), 
        .IN4(\mem[3][13] ), .S0(n1801), .S1(n1822), .Q(n1604) );
  MUX41X1 U1823 ( .IN1(n1604), .IN3(n1602), .IN2(n1603), .IN4(n1601), .S0(N18), 
        .S1(n1788), .Q(n1605) );
  MUX21X1 U1824 ( .IN1(n1605), .IN2(n1600), .S(N19), .Q(rd_dataB[13]) );
  MUX41X1 U1825 ( .IN1(\mem[28][14] ), .IN3(\mem[30][14] ), .IN2(\mem[29][14] ), .IN4(\mem[31][14] ), .S0(n1802), .S1(n1823), .Q(n1606) );
  MUX41X1 U1826 ( .IN1(\mem[24][14] ), .IN3(\mem[26][14] ), .IN2(\mem[25][14] ), .IN4(\mem[27][14] ), .S0(n1802), .S1(n1823), .Q(n1607) );
  MUX41X1 U1827 ( .IN1(\mem[20][14] ), .IN3(\mem[22][14] ), .IN2(\mem[21][14] ), .IN4(\mem[23][14] ), .S0(n1802), .S1(n1823), .Q(n1608) );
  MUX41X1 U1828 ( .IN1(\mem[16][14] ), .IN3(\mem[18][14] ), .IN2(\mem[17][14] ), .IN4(\mem[19][14] ), .S0(n1802), .S1(n1823), .Q(n1609) );
  MUX41X1 U1829 ( .IN1(n1609), .IN3(n1607), .IN2(n1608), .IN4(n1606), .S0(N18), 
        .S1(n1788), .Q(n1610) );
  MUX41X1 U1830 ( .IN1(\mem[12][14] ), .IN3(\mem[14][14] ), .IN2(\mem[13][14] ), .IN4(\mem[15][14] ), .S0(n1802), .S1(n1823), .Q(n1611) );
  MUX41X1 U1831 ( .IN1(\mem[8][14] ), .IN3(\mem[10][14] ), .IN2(\mem[9][14] ), 
        .IN4(\mem[11][14] ), .S0(n1802), .S1(n1823), .Q(n1612) );
  MUX41X1 U1832 ( .IN1(\mem[4][14] ), .IN3(\mem[6][14] ), .IN2(\mem[5][14] ), 
        .IN4(\mem[7][14] ), .S0(n1802), .S1(n1823), .Q(n1613) );
  MUX41X1 U1833 ( .IN1(\mem[0][14] ), .IN3(\mem[2][14] ), .IN2(\mem[1][14] ), 
        .IN4(\mem[3][14] ), .S0(n1802), .S1(n1823), .Q(n1614) );
  MUX41X1 U1834 ( .IN1(n1614), .IN3(n1612), .IN2(n1613), .IN4(n1611), .S0(N18), 
        .S1(n1788), .Q(n1615) );
  MUX21X1 U1835 ( .IN1(n1615), .IN2(n1610), .S(N19), .Q(rd_dataB[14]) );
  MUX41X1 U1836 ( .IN1(\mem[28][15] ), .IN3(\mem[30][15] ), .IN2(\mem[29][15] ), .IN4(\mem[31][15] ), .S0(n1802), .S1(n1823), .Q(n1616) );
  MUX41X1 U1837 ( .IN1(\mem[24][15] ), .IN3(\mem[26][15] ), .IN2(\mem[25][15] ), .IN4(\mem[27][15] ), .S0(n1802), .S1(n1823), .Q(n1617) );
  MUX41X1 U1838 ( .IN1(\mem[20][15] ), .IN3(\mem[22][15] ), .IN2(\mem[21][15] ), .IN4(\mem[23][15] ), .S0(n1802), .S1(n1823), .Q(n1618) );
  MUX41X1 U1839 ( .IN1(\mem[16][15] ), .IN3(\mem[18][15] ), .IN2(\mem[17][15] ), .IN4(\mem[19][15] ), .S0(n1802), .S1(n1823), .Q(n1619) );
  MUX41X1 U1840 ( .IN1(n1619), .IN3(n1617), .IN2(n1618), .IN4(n1616), .S0(N18), 
        .S1(n1788), .Q(n1620) );
  MUX41X1 U1841 ( .IN1(\mem[12][15] ), .IN3(\mem[14][15] ), .IN2(\mem[13][15] ), .IN4(\mem[15][15] ), .S0(n1811), .S1(n1824), .Q(n1621) );
  MUX41X1 U1842 ( .IN1(\mem[8][15] ), .IN3(\mem[10][15] ), .IN2(\mem[9][15] ), 
        .IN4(\mem[11][15] ), .S0(n1807), .S1(n1824), .Q(n1622) );
  MUX41X1 U1843 ( .IN1(\mem[4][15] ), .IN3(\mem[6][15] ), .IN2(\mem[5][15] ), 
        .IN4(\mem[7][15] ), .S0(n1795), .S1(n1824), .Q(n1623) );
  MUX41X1 U1844 ( .IN1(\mem[0][15] ), .IN3(\mem[2][15] ), .IN2(\mem[1][15] ), 
        .IN4(\mem[3][15] ), .S0(n1800), .S1(n1824), .Q(n1624) );
  MUX41X1 U1845 ( .IN1(n1624), .IN3(n1622), .IN2(n1623), .IN4(n1621), .S0(N18), 
        .S1(n1788), .Q(n1625) );
  MUX21X1 U1846 ( .IN1(n1625), .IN2(n1620), .S(N19), .Q(rd_dataB[15]) );
  MUX41X1 U1847 ( .IN1(\mem[28][16] ), .IN3(\mem[30][16] ), .IN2(\mem[29][16] ), .IN4(\mem[31][16] ), .S0(n1809), .S1(n1824), .Q(n1626) );
  MUX41X1 U1848 ( .IN1(\mem[24][16] ), .IN3(\mem[26][16] ), .IN2(\mem[25][16] ), .IN4(\mem[27][16] ), .S0(n1799), .S1(n1824), .Q(n1627) );
  MUX41X1 U1849 ( .IN1(\mem[20][16] ), .IN3(\mem[22][16] ), .IN2(\mem[21][16] ), .IN4(\mem[23][16] ), .S0(n1797), .S1(n1824), .Q(n1628) );
  MUX41X1 U1850 ( .IN1(\mem[16][16] ), .IN3(\mem[18][16] ), .IN2(\mem[17][16] ), .IN4(\mem[19][16] ), .S0(n1802), .S1(n1824), .Q(n1629) );
  MUX41X1 U1851 ( .IN1(n1629), .IN3(n1627), .IN2(n1628), .IN4(n1626), .S0(N18), 
        .S1(n1788), .Q(n1630) );
  MUX41X1 U1852 ( .IN1(\mem[12][16] ), .IN3(\mem[14][16] ), .IN2(\mem[13][16] ), .IN4(\mem[15][16] ), .S0(n1810), .S1(n1824), .Q(n1631) );
  MUX41X1 U1853 ( .IN1(\mem[8][16] ), .IN3(\mem[10][16] ), .IN2(\mem[9][16] ), 
        .IN4(\mem[11][16] ), .S0(n1803), .S1(n1824), .Q(n1632) );
  MUX41X1 U1854 ( .IN1(\mem[4][16] ), .IN3(\mem[6][16] ), .IN2(\mem[5][16] ), 
        .IN4(\mem[7][16] ), .S0(n1801), .S1(n1824), .Q(n1633) );
  MUX41X1 U1855 ( .IN1(\mem[0][16] ), .IN3(\mem[2][16] ), .IN2(\mem[1][16] ), 
        .IN4(\mem[3][16] ), .S0(n1798), .S1(n1824), .Q(n1634) );
  MUX41X1 U1856 ( .IN1(n1634), .IN3(n1632), .IN2(n1633), .IN4(n1631), .S0(N18), 
        .S1(n1788), .Q(n1635) );
  MUX21X1 U1857 ( .IN1(n1635), .IN2(n1630), .S(N19), .Q(rd_dataB[16]) );
  MUX41X1 U1858 ( .IN1(\mem[28][17] ), .IN3(\mem[30][17] ), .IN2(\mem[29][17] ), .IN4(\mem[31][17] ), .S0(n1803), .S1(n1825), .Q(n1636) );
  MUX41X1 U1859 ( .IN1(\mem[24][17] ), .IN3(\mem[26][17] ), .IN2(\mem[25][17] ), .IN4(\mem[27][17] ), .S0(n1803), .S1(n1825), .Q(n1637) );
  MUX41X1 U1860 ( .IN1(\mem[20][17] ), .IN3(\mem[22][17] ), .IN2(\mem[21][17] ), .IN4(\mem[23][17] ), .S0(n1803), .S1(n1825), .Q(n1638) );
  MUX41X1 U1861 ( .IN1(\mem[16][17] ), .IN3(\mem[18][17] ), .IN2(\mem[17][17] ), .IN4(\mem[19][17] ), .S0(n1803), .S1(n1825), .Q(n1639) );
  MUX41X1 U1862 ( .IN1(n1639), .IN3(n1637), .IN2(n1638), .IN4(n1636), .S0(N18), 
        .S1(n1788), .Q(n1640) );
  MUX41X1 U1863 ( .IN1(\mem[12][17] ), .IN3(\mem[14][17] ), .IN2(\mem[13][17] ), .IN4(\mem[15][17] ), .S0(n1803), .S1(n1825), .Q(n1641) );
  MUX41X1 U1864 ( .IN1(\mem[8][17] ), .IN3(\mem[10][17] ), .IN2(\mem[9][17] ), 
        .IN4(\mem[11][17] ), .S0(n1803), .S1(n1825), .Q(n1642) );
  MUX41X1 U1865 ( .IN1(\mem[4][17] ), .IN3(\mem[6][17] ), .IN2(\mem[5][17] ), 
        .IN4(\mem[7][17] ), .S0(n1803), .S1(n1825), .Q(n1643) );
  MUX41X1 U1866 ( .IN1(\mem[0][17] ), .IN3(\mem[2][17] ), .IN2(\mem[1][17] ), 
        .IN4(\mem[3][17] ), .S0(n1803), .S1(n1825), .Q(n1644) );
  MUX41X1 U1867 ( .IN1(n1644), .IN3(n1642), .IN2(n1643), .IN4(n1641), .S0(N18), 
        .S1(n1788), .Q(n1645) );
  MUX21X1 U1868 ( .IN1(n1645), .IN2(n1640), .S(N19), .Q(rd_dataB[17]) );
  MUX41X1 U1869 ( .IN1(\mem[28][18] ), .IN3(\mem[30][18] ), .IN2(\mem[29][18] ), .IN4(\mem[31][18] ), .S0(n1803), .S1(n1825), .Q(n1646) );
  MUX41X1 U1870 ( .IN1(\mem[24][18] ), .IN3(\mem[26][18] ), .IN2(\mem[25][18] ), .IN4(\mem[27][18] ), .S0(n1803), .S1(n1825), .Q(n1647) );
  MUX41X1 U1871 ( .IN1(\mem[20][18] ), .IN3(\mem[22][18] ), .IN2(\mem[21][18] ), .IN4(\mem[23][18] ), .S0(n1803), .S1(n1825), .Q(n1648) );
  MUX41X1 U1872 ( .IN1(\mem[16][18] ), .IN3(\mem[18][18] ), .IN2(\mem[17][18] ), .IN4(\mem[19][18] ), .S0(n1803), .S1(n1825), .Q(n1649) );
  MUX41X1 U1873 ( .IN1(n1649), .IN3(n1647), .IN2(n1648), .IN4(n1646), .S0(N18), 
        .S1(n1787), .Q(n1650) );
  MUX41X1 U1874 ( .IN1(\mem[12][18] ), .IN3(\mem[14][18] ), .IN2(\mem[13][18] ), .IN4(\mem[15][18] ), .S0(n1804), .S1(n1826), .Q(n1651) );
  MUX41X1 U1875 ( .IN1(\mem[8][18] ), .IN3(\mem[10][18] ), .IN2(\mem[9][18] ), 
        .IN4(\mem[11][18] ), .S0(n1804), .S1(n1826), .Q(n1652) );
  MUX41X1 U1876 ( .IN1(\mem[4][18] ), .IN3(\mem[6][18] ), .IN2(\mem[5][18] ), 
        .IN4(\mem[7][18] ), .S0(n1804), .S1(n1826), .Q(n1653) );
  MUX41X1 U1877 ( .IN1(\mem[0][18] ), .IN3(\mem[2][18] ), .IN2(\mem[1][18] ), 
        .IN4(\mem[3][18] ), .S0(n1804), .S1(n1826), .Q(n1654) );
  MUX41X1 U1878 ( .IN1(n1654), .IN3(n1652), .IN2(n1653), .IN4(n1651), .S0(N18), 
        .S1(n1787), .Q(n1655) );
  MUX21X1 U1879 ( .IN1(n1655), .IN2(n1650), .S(N19), .Q(rd_dataB[18]) );
  MUX41X1 U1880 ( .IN1(\mem[28][19] ), .IN3(\mem[30][19] ), .IN2(\mem[29][19] ), .IN4(\mem[31][19] ), .S0(n1804), .S1(n1826), .Q(n1656) );
  MUX41X1 U1881 ( .IN1(\mem[24][19] ), .IN3(\mem[26][19] ), .IN2(\mem[25][19] ), .IN4(\mem[27][19] ), .S0(n1804), .S1(n1826), .Q(n1657) );
  MUX41X1 U1882 ( .IN1(\mem[20][19] ), .IN3(\mem[22][19] ), .IN2(\mem[21][19] ), .IN4(\mem[23][19] ), .S0(n1804), .S1(n1826), .Q(n1658) );
  MUX41X1 U1883 ( .IN1(\mem[16][19] ), .IN3(\mem[18][19] ), .IN2(\mem[17][19] ), .IN4(\mem[19][19] ), .S0(n1804), .S1(n1826), .Q(n1659) );
  MUX41X1 U1884 ( .IN1(n1659), .IN3(n1657), .IN2(n1658), .IN4(n1656), .S0(N18), 
        .S1(n1787), .Q(n1660) );
  MUX41X1 U1885 ( .IN1(\mem[12][19] ), .IN3(\mem[14][19] ), .IN2(\mem[13][19] ), .IN4(\mem[15][19] ), .S0(n1804), .S1(n1826), .Q(n1661) );
  MUX41X1 U1886 ( .IN1(\mem[8][19] ), .IN3(\mem[10][19] ), .IN2(\mem[9][19] ), 
        .IN4(\mem[11][19] ), .S0(n1804), .S1(n1826), .Q(n1662) );
  MUX41X1 U1887 ( .IN1(\mem[4][19] ), .IN3(\mem[6][19] ), .IN2(\mem[5][19] ), 
        .IN4(\mem[7][19] ), .S0(n1804), .S1(n1826), .Q(n1663) );
  MUX41X1 U1888 ( .IN1(\mem[0][19] ), .IN3(\mem[2][19] ), .IN2(\mem[1][19] ), 
        .IN4(\mem[3][19] ), .S0(n1804), .S1(n1826), .Q(n1664) );
  MUX41X1 U1889 ( .IN1(n1664), .IN3(n1662), .IN2(n1663), .IN4(n1661), .S0(N18), 
        .S1(n1787), .Q(n1665) );
  MUX21X1 U1890 ( .IN1(n1665), .IN2(n1660), .S(N19), .Q(rd_dataB[19]) );
  MUX41X1 U1891 ( .IN1(\mem[28][20] ), .IN3(\mem[30][20] ), .IN2(\mem[29][20] ), .IN4(\mem[31][20] ), .S0(n1805), .S1(n1827), .Q(n1666) );
  MUX41X1 U1892 ( .IN1(\mem[24][20] ), .IN3(\mem[26][20] ), .IN2(\mem[25][20] ), .IN4(\mem[27][20] ), .S0(n1805), .S1(n1827), .Q(n1667) );
  MUX41X1 U1893 ( .IN1(\mem[20][20] ), .IN3(\mem[22][20] ), .IN2(\mem[21][20] ), .IN4(\mem[23][20] ), .S0(n1805), .S1(n1827), .Q(n1668) );
  MUX41X1 U1894 ( .IN1(\mem[16][20] ), .IN3(\mem[18][20] ), .IN2(\mem[17][20] ), .IN4(\mem[19][20] ), .S0(n1805), .S1(n1827), .Q(n1669) );
  MUX41X1 U1895 ( .IN1(n1669), .IN3(n1667), .IN2(n1668), .IN4(n1666), .S0(N18), 
        .S1(n1787), .Q(n1670) );
  MUX41X1 U1896 ( .IN1(\mem[12][20] ), .IN3(\mem[14][20] ), .IN2(\mem[13][20] ), .IN4(\mem[15][20] ), .S0(n1805), .S1(n1827), .Q(n1671) );
  MUX41X1 U1897 ( .IN1(\mem[8][20] ), .IN3(\mem[10][20] ), .IN2(\mem[9][20] ), 
        .IN4(\mem[11][20] ), .S0(n1805), .S1(n1827), .Q(n1672) );
  MUX41X1 U1898 ( .IN1(\mem[4][20] ), .IN3(\mem[6][20] ), .IN2(\mem[5][20] ), 
        .IN4(\mem[7][20] ), .S0(n1805), .S1(n1827), .Q(n1673) );
  MUX41X1 U1899 ( .IN1(\mem[0][20] ), .IN3(\mem[2][20] ), .IN2(\mem[1][20] ), 
        .IN4(\mem[3][20] ), .S0(n1805), .S1(n1827), .Q(n1674) );
  MUX41X1 U1900 ( .IN1(n1674), .IN3(n1672), .IN2(n1673), .IN4(n1671), .S0(N18), 
        .S1(n1787), .Q(n1675) );
  MUX21X1 U1901 ( .IN1(n1675), .IN2(n1670), .S(N19), .Q(rd_dataB[20]) );
  MUX41X1 U1902 ( .IN1(\mem[28][21] ), .IN3(\mem[30][21] ), .IN2(\mem[29][21] ), .IN4(\mem[31][21] ), .S0(n1805), .S1(n1827), .Q(n1676) );
  MUX41X1 U1903 ( .IN1(\mem[24][21] ), .IN3(\mem[26][21] ), .IN2(\mem[25][21] ), .IN4(\mem[27][21] ), .S0(n1805), .S1(n1827), .Q(n1677) );
  MUX41X1 U1904 ( .IN1(\mem[20][21] ), .IN3(\mem[22][21] ), .IN2(\mem[21][21] ), .IN4(\mem[23][21] ), .S0(n1805), .S1(n1827), .Q(n1678) );
  MUX41X1 U1905 ( .IN1(\mem[16][21] ), .IN3(\mem[18][21] ), .IN2(\mem[17][21] ), .IN4(\mem[19][21] ), .S0(n1805), .S1(n1827), .Q(n1679) );
  MUX41X1 U1906 ( .IN1(n1679), .IN3(n1677), .IN2(n1678), .IN4(n1676), .S0(N18), 
        .S1(n1787), .Q(n1680) );
  MUX41X1 U1907 ( .IN1(\mem[12][21] ), .IN3(\mem[14][21] ), .IN2(\mem[13][21] ), .IN4(\mem[15][21] ), .S0(n1806), .S1(n1828), .Q(n1681) );
  MUX41X1 U1908 ( .IN1(\mem[8][21] ), .IN3(\mem[10][21] ), .IN2(\mem[9][21] ), 
        .IN4(\mem[11][21] ), .S0(n1806), .S1(n1828), .Q(n1682) );
  MUX41X1 U1909 ( .IN1(\mem[4][21] ), .IN3(\mem[6][21] ), .IN2(\mem[5][21] ), 
        .IN4(\mem[7][21] ), .S0(n1806), .S1(n1828), .Q(n1683) );
  MUX41X1 U1910 ( .IN1(\mem[0][21] ), .IN3(\mem[2][21] ), .IN2(\mem[1][21] ), 
        .IN4(\mem[3][21] ), .S0(n1806), .S1(n1828), .Q(n1684) );
  MUX41X1 U1911 ( .IN1(n1684), .IN3(n1682), .IN2(n1683), .IN4(n1681), .S0(N18), 
        .S1(n1787), .Q(n1685) );
  MUX21X1 U1912 ( .IN1(n1685), .IN2(n1680), .S(N19), .Q(rd_dataB[21]) );
  MUX41X1 U1913 ( .IN1(\mem[28][22] ), .IN3(\mem[30][22] ), .IN2(\mem[29][22] ), .IN4(\mem[31][22] ), .S0(n1806), .S1(n1828), .Q(n1686) );
  MUX41X1 U1914 ( .IN1(\mem[24][22] ), .IN3(\mem[26][22] ), .IN2(\mem[25][22] ), .IN4(\mem[27][22] ), .S0(n1806), .S1(n1828), .Q(n1687) );
  MUX41X1 U1915 ( .IN1(\mem[20][22] ), .IN3(\mem[22][22] ), .IN2(\mem[21][22] ), .IN4(\mem[23][22] ), .S0(n1806), .S1(n1828), .Q(n1688) );
  MUX41X1 U1916 ( .IN1(\mem[16][22] ), .IN3(\mem[18][22] ), .IN2(\mem[17][22] ), .IN4(\mem[19][22] ), .S0(n1806), .S1(n1828), .Q(n1689) );
  MUX41X1 U1917 ( .IN1(n1689), .IN3(n1687), .IN2(n1688), .IN4(n1686), .S0(N18), 
        .S1(n1787), .Q(n1690) );
  MUX41X1 U1918 ( .IN1(\mem[12][22] ), .IN3(\mem[14][22] ), .IN2(\mem[13][22] ), .IN4(\mem[15][22] ), .S0(n1806), .S1(n1828), .Q(n1691) );
  MUX41X1 U1919 ( .IN1(\mem[8][22] ), .IN3(\mem[10][22] ), .IN2(\mem[9][22] ), 
        .IN4(\mem[11][22] ), .S0(n1806), .S1(n1828), .Q(n1692) );
  MUX41X1 U1920 ( .IN1(\mem[4][22] ), .IN3(\mem[6][22] ), .IN2(\mem[5][22] ), 
        .IN4(\mem[7][22] ), .S0(n1806), .S1(n1828), .Q(n1693) );
  MUX41X1 U1921 ( .IN1(\mem[0][22] ), .IN3(\mem[2][22] ), .IN2(\mem[1][22] ), 
        .IN4(\mem[3][22] ), .S0(n1806), .S1(n1828), .Q(n1694) );
  MUX41X1 U1922 ( .IN1(n1694), .IN3(n1692), .IN2(n1693), .IN4(n1691), .S0(N18), 
        .S1(n1787), .Q(n1695) );
  MUX21X1 U1923 ( .IN1(n1695), .IN2(n1690), .S(N19), .Q(rd_dataB[22]) );
  MUX41X1 U1924 ( .IN1(\mem[28][23] ), .IN3(\mem[30][23] ), .IN2(\mem[29][23] ), .IN4(\mem[31][23] ), .S0(n1807), .S1(n1829), .Q(n1696) );
  MUX41X1 U1925 ( .IN1(\mem[24][23] ), .IN3(\mem[26][23] ), .IN2(\mem[25][23] ), .IN4(\mem[27][23] ), .S0(n1807), .S1(n1829), .Q(n1697) );
  MUX41X1 U1926 ( .IN1(\mem[20][23] ), .IN3(\mem[22][23] ), .IN2(\mem[21][23] ), .IN4(\mem[23][23] ), .S0(n1807), .S1(n1829), .Q(n1698) );
  MUX41X1 U1927 ( .IN1(\mem[16][23] ), .IN3(\mem[18][23] ), .IN2(\mem[17][23] ), .IN4(\mem[19][23] ), .S0(n1807), .S1(n1829), .Q(n1699) );
  MUX41X1 U1928 ( .IN1(n1699), .IN3(n1697), .IN2(n1698), .IN4(n1696), .S0(N18), 
        .S1(n1787), .Q(n1700) );
  MUX41X1 U1929 ( .IN1(\mem[12][23] ), .IN3(\mem[14][23] ), .IN2(\mem[13][23] ), .IN4(\mem[15][23] ), .S0(n1807), .S1(n1829), .Q(n1701) );
  MUX41X1 U1930 ( .IN1(\mem[8][23] ), .IN3(\mem[10][23] ), .IN2(\mem[9][23] ), 
        .IN4(\mem[11][23] ), .S0(n1807), .S1(n1829), .Q(n1702) );
  MUX41X1 U1931 ( .IN1(\mem[4][23] ), .IN3(\mem[6][23] ), .IN2(\mem[5][23] ), 
        .IN4(\mem[7][23] ), .S0(n1807), .S1(n1829), .Q(n1703) );
  MUX41X1 U1932 ( .IN1(\mem[0][23] ), .IN3(\mem[2][23] ), .IN2(\mem[1][23] ), 
        .IN4(\mem[3][23] ), .S0(n1807), .S1(n1829), .Q(n1704) );
  MUX41X1 U1933 ( .IN1(n1704), .IN3(n1702), .IN2(n1703), .IN4(n1701), .S0(N18), 
        .S1(n1787), .Q(n1705) );
  MUX21X1 U1934 ( .IN1(n1705), .IN2(n1700), .S(N19), .Q(rd_dataB[23]) );
  MUX41X1 U1935 ( .IN1(\mem[28][24] ), .IN3(\mem[30][24] ), .IN2(\mem[29][24] ), .IN4(\mem[31][24] ), .S0(n1807), .S1(n1829), .Q(n1706) );
  MUX41X1 U1936 ( .IN1(\mem[24][24] ), .IN3(\mem[26][24] ), .IN2(\mem[25][24] ), .IN4(\mem[27][24] ), .S0(n1807), .S1(n1829), .Q(n1707) );
  MUX41X1 U1937 ( .IN1(\mem[20][24] ), .IN3(\mem[22][24] ), .IN2(\mem[21][24] ), .IN4(\mem[23][24] ), .S0(n1807), .S1(n1829), .Q(n1708) );
  MUX41X1 U1938 ( .IN1(\mem[16][24] ), .IN3(\mem[18][24] ), .IN2(\mem[17][24] ), .IN4(\mem[19][24] ), .S0(n1807), .S1(n1829), .Q(n1709) );
  MUX41X1 U1939 ( .IN1(n1709), .IN3(n1707), .IN2(n1708), .IN4(n1706), .S0(N18), 
        .S1(N17), .Q(n1710) );
  MUX41X1 U1940 ( .IN1(\mem[12][24] ), .IN3(\mem[14][24] ), .IN2(\mem[13][24] ), .IN4(\mem[15][24] ), .S0(n1808), .S1(n1830), .Q(n1711) );
  MUX41X1 U1941 ( .IN1(\mem[8][24] ), .IN3(\mem[10][24] ), .IN2(\mem[9][24] ), 
        .IN4(\mem[11][24] ), .S0(n1808), .S1(n1830), .Q(n1712) );
  MUX41X1 U1942 ( .IN1(\mem[4][24] ), .IN3(\mem[6][24] ), .IN2(\mem[5][24] ), 
        .IN4(\mem[7][24] ), .S0(n1808), .S1(n1830), .Q(n1713) );
  MUX41X1 U1943 ( .IN1(\mem[0][24] ), .IN3(\mem[2][24] ), .IN2(\mem[1][24] ), 
        .IN4(\mem[3][24] ), .S0(n1808), .S1(n1830), .Q(n1714) );
  MUX41X1 U1944 ( .IN1(n1714), .IN3(n1712), .IN2(n1713), .IN4(n1711), .S0(N18), 
        .S1(N17), .Q(n1715) );
  MUX21X1 U1945 ( .IN1(n1715), .IN2(n1710), .S(N19), .Q(rd_dataB[24]) );
  MUX41X1 U1946 ( .IN1(\mem[28][25] ), .IN3(\mem[30][25] ), .IN2(\mem[29][25] ), .IN4(\mem[31][25] ), .S0(n1808), .S1(n1830), .Q(n1716) );
  MUX41X1 U1947 ( .IN1(\mem[24][25] ), .IN3(\mem[26][25] ), .IN2(\mem[25][25] ), .IN4(\mem[27][25] ), .S0(n1808), .S1(n1830), .Q(n1717) );
  MUX41X1 U1948 ( .IN1(\mem[20][25] ), .IN3(\mem[22][25] ), .IN2(\mem[21][25] ), .IN4(\mem[23][25] ), .S0(n1808), .S1(n1830), .Q(n1718) );
  MUX41X1 U1949 ( .IN1(\mem[16][25] ), .IN3(\mem[18][25] ), .IN2(\mem[17][25] ), .IN4(\mem[19][25] ), .S0(n1808), .S1(n1830), .Q(n1719) );
  MUX41X1 U1950 ( .IN1(n1719), .IN3(n1717), .IN2(n1718), .IN4(n1716), .S0(N18), 
        .S1(N17), .Q(n1720) );
  MUX41X1 U1951 ( .IN1(\mem[12][25] ), .IN3(\mem[14][25] ), .IN2(\mem[13][25] ), .IN4(\mem[15][25] ), .S0(n1808), .S1(n1830), .Q(n1721) );
  MUX41X1 U1952 ( .IN1(\mem[8][25] ), .IN3(\mem[10][25] ), .IN2(\mem[9][25] ), 
        .IN4(\mem[11][25] ), .S0(n1808), .S1(n1830), .Q(n1722) );
  MUX41X1 U1953 ( .IN1(\mem[4][25] ), .IN3(\mem[6][25] ), .IN2(\mem[5][25] ), 
        .IN4(\mem[7][25] ), .S0(n1808), .S1(n1830), .Q(n1723) );
  MUX41X1 U1954 ( .IN1(\mem[0][25] ), .IN3(\mem[2][25] ), .IN2(\mem[1][25] ), 
        .IN4(\mem[3][25] ), .S0(n1808), .S1(n1830), .Q(n1724) );
  MUX41X1 U1955 ( .IN1(n1724), .IN3(n1722), .IN2(n1723), .IN4(n1721), .S0(N18), 
        .S1(N17), .Q(n1725) );
  MUX21X1 U1956 ( .IN1(n1725), .IN2(n1720), .S(N19), .Q(rd_dataB[25]) );
  MUX41X1 U1957 ( .IN1(\mem[28][26] ), .IN3(\mem[30][26] ), .IN2(\mem[29][26] ), .IN4(\mem[31][26] ), .S0(n1809), .S1(n1831), .Q(n1726) );
  MUX41X1 U1958 ( .IN1(\mem[24][26] ), .IN3(\mem[26][26] ), .IN2(\mem[25][26] ), .IN4(\mem[27][26] ), .S0(n1809), .S1(n1831), .Q(n1727) );
  MUX41X1 U1959 ( .IN1(\mem[20][26] ), .IN3(\mem[22][26] ), .IN2(\mem[21][26] ), .IN4(\mem[23][26] ), .S0(n1809), .S1(n1831), .Q(n1728) );
  MUX41X1 U1960 ( .IN1(\mem[16][26] ), .IN3(\mem[18][26] ), .IN2(\mem[17][26] ), .IN4(\mem[19][26] ), .S0(n1809), .S1(n1831), .Q(n1729) );
  MUX41X1 U1961 ( .IN1(n1729), .IN3(n1727), .IN2(n1728), .IN4(n1726), .S0(N18), 
        .S1(n1788), .Q(n1730) );
  MUX41X1 U1962 ( .IN1(\mem[12][26] ), .IN3(\mem[14][26] ), .IN2(\mem[13][26] ), .IN4(\mem[15][26] ), .S0(n1809), .S1(n1831), .Q(n1731) );
  MUX41X1 U1963 ( .IN1(\mem[8][26] ), .IN3(\mem[10][26] ), .IN2(\mem[9][26] ), 
        .IN4(\mem[11][26] ), .S0(n1809), .S1(n1831), .Q(n1732) );
  MUX41X1 U1964 ( .IN1(\mem[4][26] ), .IN3(\mem[6][26] ), .IN2(\mem[5][26] ), 
        .IN4(\mem[7][26] ), .S0(n1809), .S1(n1831), .Q(n1733) );
  MUX41X1 U1965 ( .IN1(\mem[0][26] ), .IN3(\mem[2][26] ), .IN2(\mem[1][26] ), 
        .IN4(\mem[3][26] ), .S0(n1809), .S1(n1831), .Q(n1734) );
  MUX41X1 U1966 ( .IN1(n1734), .IN3(n1732), .IN2(n1733), .IN4(n1731), .S0(N18), 
        .S1(N17), .Q(n1735) );
  MUX21X1 U1967 ( .IN1(n1735), .IN2(n1730), .S(N19), .Q(rd_dataB[26]) );
  MUX41X1 U1968 ( .IN1(\mem[28][27] ), .IN3(\mem[30][27] ), .IN2(\mem[29][27] ), .IN4(\mem[31][27] ), .S0(n1809), .S1(n1831), .Q(n1736) );
  MUX41X1 U1969 ( .IN1(\mem[24][27] ), .IN3(\mem[26][27] ), .IN2(\mem[25][27] ), .IN4(\mem[27][27] ), .S0(n1809), .S1(n1831), .Q(n1737) );
  MUX41X1 U1970 ( .IN1(\mem[20][27] ), .IN3(\mem[22][27] ), .IN2(\mem[21][27] ), .IN4(\mem[23][27] ), .S0(n1809), .S1(n1831), .Q(n1738) );
  MUX41X1 U1971 ( .IN1(\mem[16][27] ), .IN3(\mem[18][27] ), .IN2(\mem[17][27] ), .IN4(\mem[19][27] ), .S0(n1809), .S1(n1831), .Q(n1739) );
  MUX41X1 U1972 ( .IN1(n1739), .IN3(n1737), .IN2(n1738), .IN4(n1736), .S0(N18), 
        .S1(N17), .Q(n1740) );
  MUX41X1 U1973 ( .IN1(\mem[12][27] ), .IN3(\mem[14][27] ), .IN2(\mem[13][27] ), .IN4(\mem[15][27] ), .S0(n1810), .S1(n1832), .Q(n1741) );
  MUX41X1 U1974 ( .IN1(\mem[8][27] ), .IN3(\mem[10][27] ), .IN2(\mem[9][27] ), 
        .IN4(\mem[11][27] ), .S0(n1810), .S1(n1832), .Q(n1742) );
  MUX41X1 U1975 ( .IN1(\mem[4][27] ), .IN3(\mem[6][27] ), .IN2(\mem[5][27] ), 
        .IN4(\mem[7][27] ), .S0(n1810), .S1(n1832), .Q(n1743) );
  MUX41X1 U1976 ( .IN1(\mem[0][27] ), .IN3(\mem[2][27] ), .IN2(\mem[1][27] ), 
        .IN4(\mem[3][27] ), .S0(n1810), .S1(n1832), .Q(n1744) );
  MUX41X1 U1977 ( .IN1(n1744), .IN3(n1742), .IN2(n1743), .IN4(n1741), .S0(N18), 
        .S1(N17), .Q(n1745) );
  MUX21X1 U1978 ( .IN1(n1745), .IN2(n1740), .S(N19), .Q(rd_dataB[27]) );
  MUX41X1 U1979 ( .IN1(\mem[28][28] ), .IN3(\mem[30][28] ), .IN2(\mem[29][28] ), .IN4(\mem[31][28] ), .S0(n1810), .S1(n1832), .Q(n1746) );
  MUX41X1 U1980 ( .IN1(\mem[24][28] ), .IN3(\mem[26][28] ), .IN2(\mem[25][28] ), .IN4(\mem[27][28] ), .S0(n1810), .S1(n1832), .Q(n1747) );
  MUX41X1 U1981 ( .IN1(\mem[20][28] ), .IN3(\mem[22][28] ), .IN2(\mem[21][28] ), .IN4(\mem[23][28] ), .S0(n1810), .S1(n1832), .Q(n1748) );
  MUX41X1 U1982 ( .IN1(\mem[16][28] ), .IN3(\mem[18][28] ), .IN2(\mem[17][28] ), .IN4(\mem[19][28] ), .S0(n1810), .S1(n1832), .Q(n1749) );
  MUX41X1 U1983 ( .IN1(n1749), .IN3(n1747), .IN2(n1748), .IN4(n1746), .S0(N18), 
        .S1(n1787), .Q(n1750) );
  MUX41X1 U1984 ( .IN1(\mem[12][28] ), .IN3(\mem[14][28] ), .IN2(\mem[13][28] ), .IN4(\mem[15][28] ), .S0(n1810), .S1(n1832), .Q(n1751) );
  MUX41X1 U1985 ( .IN1(\mem[8][28] ), .IN3(\mem[10][28] ), .IN2(\mem[9][28] ), 
        .IN4(\mem[11][28] ), .S0(n1810), .S1(n1832), .Q(n1752) );
  MUX41X1 U1986 ( .IN1(\mem[4][28] ), .IN3(\mem[6][28] ), .IN2(\mem[5][28] ), 
        .IN4(\mem[7][28] ), .S0(n1810), .S1(n1832), .Q(n1753) );
  MUX41X1 U1987 ( .IN1(\mem[0][28] ), .IN3(\mem[2][28] ), .IN2(\mem[1][28] ), 
        .IN4(\mem[3][28] ), .S0(n1810), .S1(n1832), .Q(n1754) );
  MUX41X1 U1988 ( .IN1(n1754), .IN3(n1752), .IN2(n1753), .IN4(n1751), .S0(N18), 
        .S1(N17), .Q(n1755) );
  MUX21X1 U1989 ( .IN1(n1755), .IN2(n1750), .S(N19), .Q(rd_dataB[28]) );
  MUX41X1 U1990 ( .IN1(\mem[28][29] ), .IN3(\mem[30][29] ), .IN2(\mem[29][29] ), .IN4(\mem[31][29] ), .S0(n1794), .S1(n1833), .Q(n1756) );
  MUX41X1 U1991 ( .IN1(\mem[24][29] ), .IN3(\mem[26][29] ), .IN2(\mem[25][29] ), .IN4(\mem[27][29] ), .S0(n1804), .S1(n1833), .Q(n1757) );
  MUX41X1 U1992 ( .IN1(\mem[20][29] ), .IN3(\mem[22][29] ), .IN2(\mem[21][29] ), .IN4(\mem[23][29] ), .S0(n1806), .S1(n1833), .Q(n1758) );
  MUX41X1 U1993 ( .IN1(\mem[16][29] ), .IN3(\mem[18][29] ), .IN2(\mem[17][29] ), .IN4(\mem[19][29] ), .S0(n1803), .S1(n1833), .Q(n1759) );
  MUX41X1 U1994 ( .IN1(n1759), .IN3(n1757), .IN2(n1758), .IN4(n1756), .S0(N18), 
        .S1(N17), .Q(n1760) );
  MUX41X1 U1995 ( .IN1(\mem[12][29] ), .IN3(\mem[14][29] ), .IN2(\mem[13][29] ), .IN4(\mem[15][29] ), .S0(n1796), .S1(n1833), .Q(n1761) );
  MUX41X1 U1996 ( .IN1(\mem[8][29] ), .IN3(\mem[10][29] ), .IN2(\mem[9][29] ), 
        .IN4(\mem[11][29] ), .S0(n1808), .S1(n1833), .Q(n1762) );
  MUX41X1 U1997 ( .IN1(\mem[4][29] ), .IN3(\mem[6][29] ), .IN2(\mem[5][29] ), 
        .IN4(\mem[7][29] ), .S0(n1805), .S1(n1833), .Q(n1763) );
  MUX41X1 U1998 ( .IN1(\mem[0][29] ), .IN3(\mem[2][29] ), .IN2(\mem[1][29] ), 
        .IN4(\mem[3][29] ), .S0(n1804), .S1(n1833), .Q(n1764) );
  MUX41X1 U1999 ( .IN1(n1764), .IN3(n1762), .IN2(n1763), .IN4(n1761), .S0(N18), 
        .S1(N17), .Q(n1765) );
  MUX21X1 U2000 ( .IN1(n1765), .IN2(n1760), .S(N19), .Q(rd_dataB[29]) );
  MUX41X1 U2001 ( .IN1(\mem[28][30] ), .IN3(\mem[30][30] ), .IN2(\mem[29][30] ), .IN4(\mem[31][30] ), .S0(n1793), .S1(n1833), .Q(n1766) );
  MUX41X1 U2002 ( .IN1(\mem[24][30] ), .IN3(\mem[26][30] ), .IN2(\mem[25][30] ), .IN4(\mem[27][30] ), .S0(n1806), .S1(n1833), .Q(n1767) );
  MUX41X1 U2003 ( .IN1(\mem[20][30] ), .IN3(\mem[22][30] ), .IN2(\mem[21][30] ), .IN4(\mem[23][30] ), .S0(n1805), .S1(n1833), .Q(n1768) );
  MUX41X1 U2004 ( .IN1(\mem[16][30] ), .IN3(\mem[18][30] ), .IN2(\mem[17][30] ), .IN4(\mem[19][30] ), .S0(n1808), .S1(n1833), .Q(n1769) );
  MUX41X1 U2005 ( .IN1(n1769), .IN3(n1767), .IN2(n1768), .IN4(n1766), .S0(N18), 
        .S1(n1790), .Q(n1770) );
  MUX41X1 U2006 ( .IN1(\mem[12][30] ), .IN3(\mem[14][30] ), .IN2(\mem[13][30] ), .IN4(\mem[15][30] ), .S0(n1811), .S1(n1830), .Q(n1771) );
  MUX41X1 U2007 ( .IN1(\mem[8][30] ), .IN3(\mem[10][30] ), .IN2(\mem[9][30] ), 
        .IN4(\mem[11][30] ), .S0(n1811), .S1(n1829), .Q(n1772) );
  MUX41X1 U2008 ( .IN1(\mem[4][30] ), .IN3(\mem[6][30] ), .IN2(\mem[5][30] ), 
        .IN4(\mem[7][30] ), .S0(n1811), .S1(n1814), .Q(n1773) );
  MUX41X1 U2009 ( .IN1(\mem[0][30] ), .IN3(\mem[2][30] ), .IN2(\mem[1][30] ), 
        .IN4(\mem[3][30] ), .S0(n1811), .S1(n1828), .Q(n1774) );
  MUX41X1 U2010 ( .IN1(n1774), .IN3(n1772), .IN2(n1773), .IN4(n1771), .S0(N18), 
        .S1(N17), .Q(n1775) );
  MUX21X1 U2011 ( .IN1(n1775), .IN2(n1770), .S(N19), .Q(rd_dataB[30]) );
  MUX41X1 U2012 ( .IN1(\mem[28][31] ), .IN3(\mem[30][31] ), .IN2(\mem[29][31] ), .IN4(\mem[31][31] ), .S0(n1811), .S1(n1832), .Q(n1776) );
  MUX41X1 U2013 ( .IN1(\mem[24][31] ), .IN3(\mem[26][31] ), .IN2(\mem[25][31] ), .IN4(\mem[27][31] ), .S0(n1811), .S1(n1817), .Q(n1777) );
  MUX41X1 U2014 ( .IN1(\mem[20][31] ), .IN3(\mem[22][31] ), .IN2(\mem[21][31] ), .IN4(\mem[23][31] ), .S0(n1811), .S1(n1827), .Q(n1778) );
  MUX41X1 U2015 ( .IN1(\mem[16][31] ), .IN3(\mem[18][31] ), .IN2(\mem[17][31] ), .IN4(\mem[19][31] ), .S0(n1811), .S1(n1825), .Q(n1779) );
  MUX41X1 U2016 ( .IN1(n1779), .IN3(n1777), .IN2(n1778), .IN4(n1776), .S0(N18), 
        .S1(n1789), .Q(n1780) );
  MUX41X1 U2017 ( .IN1(\mem[12][31] ), .IN3(\mem[14][31] ), .IN2(\mem[13][31] ), .IN4(\mem[15][31] ), .S0(n1811), .S1(n1833), .Q(n1781) );
  MUX41X1 U2018 ( .IN1(\mem[8][31] ), .IN3(\mem[10][31] ), .IN2(\mem[9][31] ), 
        .IN4(\mem[11][31] ), .S0(n1811), .S1(n1831), .Q(n1782) );
  MUX41X1 U2019 ( .IN1(\mem[4][31] ), .IN3(\mem[6][31] ), .IN2(\mem[5][31] ), 
        .IN4(\mem[7][31] ), .S0(n1811), .S1(n1815), .Q(n1783) );
  MUX41X1 U2020 ( .IN1(\mem[0][31] ), .IN3(\mem[2][31] ), .IN2(\mem[1][31] ), 
        .IN4(\mem[3][31] ), .S0(n1811), .S1(n1826), .Q(n1784) );
  MUX41X1 U2021 ( .IN1(n1784), .IN3(n1782), .IN2(n1783), .IN4(n1781), .S0(N18), 
        .S1(N17), .Q(n1785) );
  MUX21X1 U2022 ( .IN1(n1785), .IN2(n1780), .S(N19), .Q(rd_dataB[31]) );
  AO21X1 U2023 ( .IN1(n86), .IN2(n73), .IN3(n1999), .Q(n1841) );
  AO21X1 U2024 ( .IN1(n86), .IN2(n73), .IN3(n1999), .Q(n1842) );
  AO21X1 U2025 ( .IN1(n83), .IN2(n73), .IN3(n1999), .Q(n1846) );
  AO21X1 U2026 ( .IN1(n83), .IN2(n73), .IN3(n1999), .Q(n1847) );
  AND2X1 U2027 ( .IN1(wr_data[23]), .IN2(n1839), .Q(n1855) );
  AND2X1 U2028 ( .IN1(wr_data[23]), .IN2(n1838), .Q(n1856) );
  AND2X1 U2029 ( .IN1(wr_data[22]), .IN2(n1836), .Q(n1857) );
  AND2X1 U2030 ( .IN1(wr_data[22]), .IN2(n1838), .Q(n1858) );
  AND2X1 U2031 ( .IN1(wr_data[21]), .IN2(n1840), .Q(n1859) );
  AND2X1 U2032 ( .IN1(wr_data[21]), .IN2(n1840), .Q(n1860) );
  AND2X1 U2033 ( .IN1(wr_data[20]), .IN2(n1834), .Q(n1861) );
  AND2X1 U2034 ( .IN1(wr_data[20]), .IN2(n1840), .Q(n1862) );
  AND2X1 U2035 ( .IN1(wr_data[19]), .IN2(n1840), .Q(n1863) );
  AND2X1 U2036 ( .IN1(wr_data[19]), .IN2(n1840), .Q(n1864) );
  AND2X1 U2037 ( .IN1(wr_data[18]), .IN2(n1834), .Q(n1865) );
  AND2X1 U2038 ( .IN1(wr_data[18]), .IN2(n1840), .Q(n1866) );
  AND2X1 U2039 ( .IN1(wr_data[17]), .IN2(n1840), .Q(n1867) );
  AND2X1 U2040 ( .IN1(wr_data[17]), .IN2(n1837), .Q(n1868) );
  AND2X1 U2041 ( .IN1(wr_data[16]), .IN2(n1834), .Q(n1869) );
  AND2X1 U2042 ( .IN1(wr_data[16]), .IN2(n1834), .Q(n1870) );
  AND2X1 U2043 ( .IN1(wr_data[15]), .IN2(n1835), .Q(n1871) );
  AND2X1 U2044 ( .IN1(wr_data[14]), .IN2(n1840), .Q(n1873) );
  AO21X1 U2045 ( .IN1(n94), .IN2(n73), .IN3(n1999), .Q(n1877) );
  AO21X1 U2046 ( .IN1(n94), .IN2(n73), .IN3(n1999), .Q(n1878) );
  AO21X1 U2047 ( .IN1(n104), .IN2(n81), .IN3(n1999), .Q(n1879) );
  AO21X1 U2048 ( .IN1(n104), .IN2(n81), .IN3(n1999), .Q(n1880) );
  AO21X1 U2049 ( .IN1(n104), .IN2(n79), .IN3(n1999), .Q(n1881) );
  AO21X1 U2050 ( .IN1(n104), .IN2(n79), .IN3(n1999), .Q(n1882) );
  AO21X1 U2051 ( .IN1(n104), .IN2(n77), .IN3(n1999), .Q(n1883) );
  AO21X1 U2052 ( .IN1(n104), .IN2(n77), .IN3(n1999), .Q(n1884) );
  AO21X1 U2053 ( .IN1(n104), .IN2(n75), .IN3(n1999), .Q(n1885) );
  AO21X1 U2054 ( .IN1(n104), .IN2(n75), .IN3(n1999), .Q(n1886) );
  AO21X1 U2055 ( .IN1(n95), .IN2(n81), .IN3(n1998), .Q(n1895) );
  AO21X1 U2056 ( .IN1(n95), .IN2(n81), .IN3(n1998), .Q(n1896) );
  AO21X1 U2057 ( .IN1(n95), .IN2(n79), .IN3(n1998), .Q(n1897) );
  AO21X1 U2058 ( .IN1(n95), .IN2(n79), .IN3(n1998), .Q(n1898) );
  AO21X1 U2059 ( .IN1(n95), .IN2(n77), .IN3(n1998), .Q(n1899) );
  AO21X1 U2060 ( .IN1(n95), .IN2(n77), .IN3(n1998), .Q(n1900) );
  AO21X1 U2061 ( .IN1(n95), .IN2(n75), .IN3(n1998), .Q(n1901) );
  AO21X1 U2062 ( .IN1(n95), .IN2(n75), .IN3(n1998), .Q(n1902) );
  AO21X1 U2063 ( .IN1(n84), .IN2(n81), .IN3(n1997), .Q(n1911) );
  AO21X1 U2064 ( .IN1(n84), .IN2(n81), .IN3(n1997), .Q(n1912) );
  AO21X1 U2065 ( .IN1(n84), .IN2(n79), .IN3(n1997), .Q(n1913) );
  AO21X1 U2066 ( .IN1(n84), .IN2(n79), .IN3(n1997), .Q(n1914) );
  AO21X1 U2067 ( .IN1(n84), .IN2(n77), .IN3(n1997), .Q(n1915) );
  AO21X1 U2068 ( .IN1(n84), .IN2(n77), .IN3(n1997), .Q(n1916) );
  AO21X1 U2069 ( .IN1(n81), .IN2(n73), .IN3(n1997), .Q(n1925) );
  AO21X1 U2070 ( .IN1(n81), .IN2(n73), .IN3(n1997), .Q(n1926) );
endmodule


module id_exe_reg ( clk, nrst, en, flush, cur_pc0, next_pc0, bra_off0, opA0, 
        opB0, mem_data0, reg_addr0, cur_pc, next_pc, bra_off, opA, opB, 
        mem_data, reg_addr );
  input [31:0] cur_pc0;
  input [31:0] next_pc0;
  input [31:0] bra_off0;
  input [31:0] opA0;
  input [31:0] opB0;
  input [31:0] mem_data0;
  input [4:0] reg_addr0;
  output [31:0] cur_pc;
  output [31:0] next_pc;
  output [31:0] bra_off;
  output [31:0] opA;
  output [31:0] opB;
  output [31:0] mem_data;
  output [4:0] reg_addr;
  input clk, nrst, en, flush;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, n2,
         n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  DFFX1 \reg_addr_reg[4]  ( .D(N199), .CLK(clk), .Q(reg_addr[4]) );
  DFFX1 \reg_addr_reg[3]  ( .D(N198), .CLK(clk), .Q(reg_addr[3]) );
  DFFX1 \reg_addr_reg[2]  ( .D(N197), .CLK(clk), .Q(reg_addr[2]) );
  DFFX1 \reg_addr_reg[1]  ( .D(N196), .CLK(clk), .Q(reg_addr[1]) );
  DFFX1 \reg_addr_reg[0]  ( .D(N195), .CLK(clk), .Q(reg_addr[0]) );
  DFFX1 \cur_pc_reg[31]  ( .D(N34), .CLK(clk), .Q(cur_pc[31]) );
  DFFX1 \cur_pc_reg[30]  ( .D(N33), .CLK(clk), .Q(cur_pc[30]) );
  DFFX1 \cur_pc_reg[29]  ( .D(N32), .CLK(clk), .Q(cur_pc[29]) );
  DFFX1 \cur_pc_reg[28]  ( .D(N31), .CLK(clk), .Q(cur_pc[28]) );
  DFFX1 \cur_pc_reg[27]  ( .D(N30), .CLK(clk), .Q(cur_pc[27]) );
  DFFX1 \cur_pc_reg[26]  ( .D(N29), .CLK(clk), .Q(cur_pc[26]) );
  DFFX1 \cur_pc_reg[25]  ( .D(N28), .CLK(clk), .Q(cur_pc[25]) );
  DFFX1 \cur_pc_reg[24]  ( .D(N27), .CLK(clk), .Q(cur_pc[24]) );
  DFFX1 \cur_pc_reg[23]  ( .D(N26), .CLK(clk), .Q(cur_pc[23]) );
  DFFX1 \cur_pc_reg[22]  ( .D(N25), .CLK(clk), .Q(cur_pc[22]) );
  DFFX1 \cur_pc_reg[21]  ( .D(N24), .CLK(clk), .Q(cur_pc[21]) );
  DFFX1 \cur_pc_reg[20]  ( .D(N23), .CLK(clk), .Q(cur_pc[20]) );
  DFFX1 \cur_pc_reg[19]  ( .D(N22), .CLK(clk), .Q(cur_pc[19]) );
  DFFX1 \cur_pc_reg[18]  ( .D(N21), .CLK(clk), .Q(cur_pc[18]) );
  DFFX1 \cur_pc_reg[17]  ( .D(N20), .CLK(clk), .Q(cur_pc[17]) );
  DFFX1 \cur_pc_reg[16]  ( .D(N19), .CLK(clk), .Q(cur_pc[16]) );
  DFFX1 \cur_pc_reg[15]  ( .D(N18), .CLK(clk), .Q(cur_pc[15]) );
  DFFX1 \cur_pc_reg[14]  ( .D(N17), .CLK(clk), .Q(cur_pc[14]) );
  DFFX1 \cur_pc_reg[13]  ( .D(N16), .CLK(clk), .Q(cur_pc[13]) );
  DFFX1 \cur_pc_reg[12]  ( .D(N15), .CLK(clk), .Q(cur_pc[12]) );
  DFFX1 \cur_pc_reg[11]  ( .D(N14), .CLK(clk), .Q(cur_pc[11]) );
  DFFX1 \cur_pc_reg[10]  ( .D(N13), .CLK(clk), .Q(cur_pc[10]) );
  DFFX1 \cur_pc_reg[9]  ( .D(N12), .CLK(clk), .Q(cur_pc[9]) );
  DFFX1 \cur_pc_reg[8]  ( .D(N11), .CLK(clk), .Q(cur_pc[8]) );
  DFFX1 \cur_pc_reg[7]  ( .D(N10), .CLK(clk), .Q(cur_pc[7]) );
  DFFX1 \cur_pc_reg[6]  ( .D(N9), .CLK(clk), .Q(cur_pc[6]) );
  DFFX1 \cur_pc_reg[5]  ( .D(N8), .CLK(clk), .Q(cur_pc[5]) );
  DFFX1 \cur_pc_reg[4]  ( .D(N7), .CLK(clk), .Q(cur_pc[4]) );
  DFFX1 \cur_pc_reg[3]  ( .D(N6), .CLK(clk), .Q(cur_pc[3]) );
  DFFX1 \cur_pc_reg[2]  ( .D(N5), .CLK(clk), .Q(cur_pc[2]) );
  DFFX1 \cur_pc_reg[1]  ( .D(N4), .CLK(clk), .Q(cur_pc[1]) );
  DFFX1 \cur_pc_reg[0]  ( .D(N3), .CLK(clk), .Q(cur_pc[0]) );
  DFFX1 \next_pc_reg[31]  ( .D(N66), .CLK(clk), .Q(next_pc[31]) );
  DFFX1 \next_pc_reg[30]  ( .D(N65), .CLK(clk), .Q(next_pc[30]) );
  DFFX1 \next_pc_reg[29]  ( .D(N64), .CLK(clk), .Q(next_pc[29]) );
  DFFX1 \next_pc_reg[28]  ( .D(N63), .CLK(clk), .Q(next_pc[28]) );
  DFFX1 \next_pc_reg[27]  ( .D(N62), .CLK(clk), .Q(next_pc[27]) );
  DFFX1 \next_pc_reg[26]  ( .D(N61), .CLK(clk), .Q(next_pc[26]) );
  DFFX1 \next_pc_reg[25]  ( .D(N60), .CLK(clk), .Q(next_pc[25]) );
  DFFX1 \next_pc_reg[24]  ( .D(N59), .CLK(clk), .Q(next_pc[24]) );
  DFFX1 \next_pc_reg[23]  ( .D(N58), .CLK(clk), .Q(next_pc[23]) );
  DFFX1 \next_pc_reg[22]  ( .D(N57), .CLK(clk), .Q(next_pc[22]) );
  DFFX1 \next_pc_reg[21]  ( .D(N56), .CLK(clk), .Q(next_pc[21]) );
  DFFX1 \next_pc_reg[20]  ( .D(N55), .CLK(clk), .Q(next_pc[20]) );
  DFFX1 \next_pc_reg[19]  ( .D(N54), .CLK(clk), .Q(next_pc[19]) );
  DFFX1 \next_pc_reg[18]  ( .D(N53), .CLK(clk), .Q(next_pc[18]) );
  DFFX1 \next_pc_reg[17]  ( .D(N52), .CLK(clk), .Q(next_pc[17]) );
  DFFX1 \next_pc_reg[16]  ( .D(N51), .CLK(clk), .Q(next_pc[16]) );
  DFFX1 \next_pc_reg[15]  ( .D(N50), .CLK(clk), .Q(next_pc[15]) );
  DFFX1 \next_pc_reg[14]  ( .D(N49), .CLK(clk), .Q(next_pc[14]) );
  DFFX1 \next_pc_reg[13]  ( .D(N48), .CLK(clk), .Q(next_pc[13]) );
  DFFX1 \next_pc_reg[12]  ( .D(N47), .CLK(clk), .Q(next_pc[12]) );
  DFFX1 \next_pc_reg[11]  ( .D(N46), .CLK(clk), .Q(next_pc[11]) );
  DFFX1 \next_pc_reg[10]  ( .D(N45), .CLK(clk), .Q(next_pc[10]) );
  DFFX1 \next_pc_reg[9]  ( .D(N44), .CLK(clk), .Q(next_pc[9]) );
  DFFX1 \next_pc_reg[8]  ( .D(N43), .CLK(clk), .Q(next_pc[8]) );
  DFFX1 \next_pc_reg[7]  ( .D(N42), .CLK(clk), .Q(next_pc[7]) );
  DFFX1 \next_pc_reg[6]  ( .D(N41), .CLK(clk), .Q(next_pc[6]) );
  DFFX1 \next_pc_reg[5]  ( .D(N40), .CLK(clk), .Q(next_pc[5]) );
  DFFX1 \next_pc_reg[4]  ( .D(N39), .CLK(clk), .Q(next_pc[4]) );
  DFFX1 \next_pc_reg[3]  ( .D(N38), .CLK(clk), .Q(next_pc[3]) );
  DFFX1 \next_pc_reg[2]  ( .D(N37), .CLK(clk), .Q(next_pc[2]) );
  DFFX1 \next_pc_reg[1]  ( .D(N36), .CLK(clk), .Q(next_pc[1]) );
  DFFX1 \next_pc_reg[0]  ( .D(N35), .CLK(clk), .Q(next_pc[0]) );
  DFFX1 \bra_off_reg[31]  ( .D(N98), .CLK(clk), .Q(bra_off[31]) );
  DFFX1 \bra_off_reg[30]  ( .D(N97), .CLK(clk), .Q(bra_off[30]) );
  DFFX1 \bra_off_reg[29]  ( .D(N96), .CLK(clk), .Q(bra_off[29]) );
  DFFX1 \bra_off_reg[28]  ( .D(N95), .CLK(clk), .Q(bra_off[28]) );
  DFFX1 \bra_off_reg[27]  ( .D(N94), .CLK(clk), .Q(bra_off[27]) );
  DFFX1 \bra_off_reg[26]  ( .D(N93), .CLK(clk), .Q(bra_off[26]) );
  DFFX1 \bra_off_reg[25]  ( .D(N92), .CLK(clk), .Q(bra_off[25]) );
  DFFX1 \bra_off_reg[24]  ( .D(N91), .CLK(clk), .Q(bra_off[24]) );
  DFFX1 \bra_off_reg[23]  ( .D(N90), .CLK(clk), .Q(bra_off[23]) );
  DFFX1 \bra_off_reg[22]  ( .D(N89), .CLK(clk), .Q(bra_off[22]) );
  DFFX1 \bra_off_reg[21]  ( .D(N88), .CLK(clk), .Q(bra_off[21]) );
  DFFX1 \bra_off_reg[20]  ( .D(N87), .CLK(clk), .Q(bra_off[20]) );
  DFFX1 \bra_off_reg[19]  ( .D(N86), .CLK(clk), .Q(bra_off[19]) );
  DFFX1 \bra_off_reg[18]  ( .D(N85), .CLK(clk), .Q(bra_off[18]) );
  DFFX1 \bra_off_reg[17]  ( .D(N84), .CLK(clk), .Q(bra_off[17]) );
  DFFX1 \bra_off_reg[16]  ( .D(N83), .CLK(clk), .Q(bra_off[16]) );
  DFFX1 \bra_off_reg[15]  ( .D(N82), .CLK(clk), .Q(bra_off[15]) );
  DFFX1 \bra_off_reg[14]  ( .D(N81), .CLK(clk), .Q(bra_off[14]) );
  DFFX1 \bra_off_reg[13]  ( .D(N80), .CLK(clk), .Q(bra_off[13]) );
  DFFX1 \bra_off_reg[12]  ( .D(N79), .CLK(clk), .Q(bra_off[12]) );
  DFFX1 \bra_off_reg[11]  ( .D(N78), .CLK(clk), .Q(bra_off[11]) );
  DFFX1 \bra_off_reg[10]  ( .D(N77), .CLK(clk), .Q(bra_off[10]) );
  DFFX1 \bra_off_reg[9]  ( .D(N76), .CLK(clk), .Q(bra_off[9]) );
  DFFX1 \bra_off_reg[8]  ( .D(N75), .CLK(clk), .Q(bra_off[8]) );
  DFFX1 \bra_off_reg[7]  ( .D(N74), .CLK(clk), .Q(bra_off[7]) );
  DFFX1 \bra_off_reg[6]  ( .D(N73), .CLK(clk), .Q(bra_off[6]) );
  DFFX1 \bra_off_reg[5]  ( .D(N72), .CLK(clk), .Q(bra_off[5]) );
  DFFX1 \bra_off_reg[4]  ( .D(N71), .CLK(clk), .Q(bra_off[4]) );
  DFFX1 \bra_off_reg[3]  ( .D(N70), .CLK(clk), .Q(bra_off[3]) );
  DFFX1 \bra_off_reg[2]  ( .D(N69), .CLK(clk), .Q(bra_off[2]) );
  DFFX1 \bra_off_reg[1]  ( .D(N68), .CLK(clk), .Q(bra_off[1]) );
  DFFX1 \bra_off_reg[0]  ( .D(N67), .CLK(clk), .Q(bra_off[0]) );
  DFFX1 \opA_reg[31]  ( .D(N130), .CLK(clk), .Q(opA[31]) );
  DFFX1 \opA_reg[30]  ( .D(N129), .CLK(clk), .Q(opA[30]) );
  DFFX1 \opA_reg[29]  ( .D(N128), .CLK(clk), .Q(opA[29]) );
  DFFX1 \opA_reg[28]  ( .D(N127), .CLK(clk), .Q(opA[28]) );
  DFFX1 \opA_reg[27]  ( .D(N126), .CLK(clk), .Q(opA[27]) );
  DFFX1 \opA_reg[26]  ( .D(N125), .CLK(clk), .Q(opA[26]) );
  DFFX1 \opA_reg[25]  ( .D(N124), .CLK(clk), .Q(opA[25]) );
  DFFX1 \opA_reg[24]  ( .D(N123), .CLK(clk), .Q(opA[24]) );
  DFFX1 \opA_reg[23]  ( .D(N122), .CLK(clk), .Q(opA[23]) );
  DFFX1 \opA_reg[22]  ( .D(N121), .CLK(clk), .Q(opA[22]) );
  DFFX1 \opA_reg[21]  ( .D(N120), .CLK(clk), .Q(opA[21]) );
  DFFX1 \opA_reg[20]  ( .D(N119), .CLK(clk), .Q(opA[20]) );
  DFFX1 \opA_reg[19]  ( .D(N118), .CLK(clk), .Q(opA[19]) );
  DFFX1 \opA_reg[18]  ( .D(N117), .CLK(clk), .Q(opA[18]) );
  DFFX1 \opA_reg[17]  ( .D(N116), .CLK(clk), .Q(opA[17]) );
  DFFX1 \opA_reg[16]  ( .D(N115), .CLK(clk), .Q(opA[16]) );
  DFFX1 \opA_reg[15]  ( .D(N114), .CLK(clk), .Q(opA[15]) );
  DFFX1 \opA_reg[14]  ( .D(N113), .CLK(clk), .Q(opA[14]) );
  DFFX1 \opA_reg[13]  ( .D(N112), .CLK(clk), .Q(opA[13]) );
  DFFX1 \opA_reg[12]  ( .D(N111), .CLK(clk), .Q(opA[12]) );
  DFFX1 \opA_reg[11]  ( .D(N110), .CLK(clk), .Q(opA[11]) );
  DFFX1 \opA_reg[10]  ( .D(N109), .CLK(clk), .Q(opA[10]) );
  DFFX1 \opA_reg[9]  ( .D(N108), .CLK(clk), .Q(opA[9]) );
  DFFX1 \opA_reg[8]  ( .D(N107), .CLK(clk), .Q(opA[8]) );
  DFFX1 \opA_reg[7]  ( .D(N106), .CLK(clk), .Q(opA[7]) );
  DFFX1 \opA_reg[6]  ( .D(N105), .CLK(clk), .Q(opA[6]) );
  DFFX1 \opA_reg[5]  ( .D(N104), .CLK(clk), .Q(opA[5]) );
  DFFX1 \opA_reg[4]  ( .D(N103), .CLK(clk), .Q(opA[4]) );
  DFFX1 \opA_reg[3]  ( .D(N102), .CLK(clk), .Q(opA[3]) );
  DFFX1 \opA_reg[2]  ( .D(N101), .CLK(clk), .Q(opA[2]) );
  DFFX1 \opA_reg[1]  ( .D(N100), .CLK(clk), .Q(opA[1]) );
  DFFX1 \opA_reg[0]  ( .D(N99), .CLK(clk), .Q(opA[0]) );
  DFFX1 \opB_reg[31]  ( .D(N162), .CLK(clk), .Q(opB[31]) );
  DFFX1 \opB_reg[30]  ( .D(N161), .CLK(clk), .Q(opB[30]) );
  DFFX1 \opB_reg[29]  ( .D(N160), .CLK(clk), .Q(opB[29]) );
  DFFX1 \opB_reg[28]  ( .D(N159), .CLK(clk), .Q(opB[28]) );
  DFFX1 \opB_reg[27]  ( .D(N158), .CLK(clk), .Q(opB[27]) );
  DFFX1 \opB_reg[26]  ( .D(N157), .CLK(clk), .Q(opB[26]) );
  DFFX1 \opB_reg[25]  ( .D(N156), .CLK(clk), .Q(opB[25]) );
  DFFX1 \opB_reg[24]  ( .D(N155), .CLK(clk), .Q(opB[24]) );
  DFFX1 \opB_reg[23]  ( .D(N154), .CLK(clk), .Q(opB[23]) );
  DFFX1 \opB_reg[22]  ( .D(N153), .CLK(clk), .Q(opB[22]) );
  DFFX1 \opB_reg[21]  ( .D(N152), .CLK(clk), .Q(opB[21]) );
  DFFX1 \opB_reg[20]  ( .D(N151), .CLK(clk), .Q(opB[20]) );
  DFFX1 \opB_reg[19]  ( .D(N150), .CLK(clk), .Q(opB[19]) );
  DFFX1 \opB_reg[18]  ( .D(N149), .CLK(clk), .Q(opB[18]) );
  DFFX1 \opB_reg[17]  ( .D(N148), .CLK(clk), .Q(opB[17]) );
  DFFX1 \opB_reg[16]  ( .D(N147), .CLK(clk), .Q(opB[16]) );
  DFFX1 \opB_reg[15]  ( .D(N146), .CLK(clk), .Q(opB[15]) );
  DFFX1 \opB_reg[14]  ( .D(N145), .CLK(clk), .Q(opB[14]) );
  DFFX1 \opB_reg[13]  ( .D(N144), .CLK(clk), .Q(opB[13]) );
  DFFX1 \opB_reg[12]  ( .D(N143), .CLK(clk), .Q(opB[12]) );
  DFFX1 \opB_reg[11]  ( .D(N142), .CLK(clk), .Q(opB[11]) );
  DFFX1 \opB_reg[10]  ( .D(N141), .CLK(clk), .Q(opB[10]) );
  DFFX1 \opB_reg[9]  ( .D(N140), .CLK(clk), .Q(opB[9]) );
  DFFX1 \opB_reg[8]  ( .D(N139), .CLK(clk), .Q(opB[8]) );
  DFFX1 \opB_reg[7]  ( .D(N138), .CLK(clk), .Q(opB[7]) );
  DFFX1 \opB_reg[6]  ( .D(N137), .CLK(clk), .Q(opB[6]) );
  DFFX1 \opB_reg[5]  ( .D(N136), .CLK(clk), .Q(opB[5]) );
  DFFX1 \opB_reg[4]  ( .D(N135), .CLK(clk), .Q(opB[4]) );
  DFFX1 \opB_reg[3]  ( .D(N134), .CLK(clk), .Q(opB[3]) );
  DFFX1 \opB_reg[2]  ( .D(N133), .CLK(clk), .Q(opB[2]) );
  DFFX1 \opB_reg[1]  ( .D(N132), .CLK(clk), .Q(opB[1]) );
  DFFX1 \opB_reg[0]  ( .D(N131), .CLK(clk), .Q(opB[0]) );
  DFFX1 \mem_data_reg[31]  ( .D(N194), .CLK(clk), .Q(mem_data[31]) );
  DFFX1 \mem_data_reg[30]  ( .D(N193), .CLK(clk), .Q(mem_data[30]) );
  DFFX1 \mem_data_reg[29]  ( .D(N192), .CLK(clk), .Q(mem_data[29]) );
  DFFX1 \mem_data_reg[28]  ( .D(N191), .CLK(clk), .Q(mem_data[28]) );
  DFFX1 \mem_data_reg[27]  ( .D(N190), .CLK(clk), .Q(mem_data[27]) );
  DFFX1 \mem_data_reg[26]  ( .D(N189), .CLK(clk), .Q(mem_data[26]) );
  DFFX1 \mem_data_reg[25]  ( .D(N188), .CLK(clk), .Q(mem_data[25]) );
  DFFX1 \mem_data_reg[24]  ( .D(N187), .CLK(clk), .Q(mem_data[24]) );
  DFFX1 \mem_data_reg[23]  ( .D(N186), .CLK(clk), .Q(mem_data[23]) );
  DFFX1 \mem_data_reg[22]  ( .D(N185), .CLK(clk), .Q(mem_data[22]) );
  DFFX1 \mem_data_reg[21]  ( .D(N184), .CLK(clk), .Q(mem_data[21]) );
  DFFX1 \mem_data_reg[20]  ( .D(N183), .CLK(clk), .Q(mem_data[20]) );
  DFFX1 \mem_data_reg[19]  ( .D(N182), .CLK(clk), .Q(mem_data[19]) );
  DFFX1 \mem_data_reg[18]  ( .D(N181), .CLK(clk), .Q(mem_data[18]) );
  DFFX1 \mem_data_reg[17]  ( .D(N180), .CLK(clk), .Q(mem_data[17]) );
  DFFX1 \mem_data_reg[16]  ( .D(N179), .CLK(clk), .Q(mem_data[16]) );
  DFFX1 \mem_data_reg[15]  ( .D(N178), .CLK(clk), .Q(mem_data[15]) );
  DFFX1 \mem_data_reg[14]  ( .D(N177), .CLK(clk), .Q(mem_data[14]) );
  DFFX1 \mem_data_reg[13]  ( .D(N176), .CLK(clk), .Q(mem_data[13]) );
  DFFX1 \mem_data_reg[12]  ( .D(N175), .CLK(clk), .Q(mem_data[12]) );
  DFFX1 \mem_data_reg[11]  ( .D(N174), .CLK(clk), .Q(mem_data[11]) );
  DFFX1 \mem_data_reg[10]  ( .D(N173), .CLK(clk), .Q(mem_data[10]) );
  DFFX1 \mem_data_reg[9]  ( .D(N172), .CLK(clk), .Q(mem_data[9]) );
  DFFX1 \mem_data_reg[8]  ( .D(N171), .CLK(clk), .Q(mem_data[8]) );
  DFFX1 \mem_data_reg[7]  ( .D(N170), .CLK(clk), .Q(mem_data[7]) );
  DFFX1 \mem_data_reg[6]  ( .D(N169), .CLK(clk), .Q(mem_data[6]) );
  DFFX1 \mem_data_reg[5]  ( .D(N168), .CLK(clk), .Q(mem_data[5]) );
  DFFX1 \mem_data_reg[4]  ( .D(N167), .CLK(clk), .Q(mem_data[4]) );
  DFFX1 \mem_data_reg[3]  ( .D(N166), .CLK(clk), .Q(mem_data[3]) );
  DFFX1 \mem_data_reg[2]  ( .D(N165), .CLK(clk), .Q(mem_data[2]) );
  DFFX1 \mem_data_reg[1]  ( .D(N164), .CLK(clk), .Q(mem_data[1]) );
  DFFX1 \mem_data_reg[0]  ( .D(N163), .CLK(clk), .Q(mem_data[0]) );
  AND2X1 U4 ( .IN1(opA0[0]), .IN2(n2), .Q(N99) );
  AND2X1 U5 ( .IN1(bra_off0[31]), .IN2(n2), .Q(N98) );
  AND2X1 U6 ( .IN1(bra_off0[30]), .IN2(n2), .Q(N97) );
  AND2X1 U7 ( .IN1(bra_off0[29]), .IN2(n2), .Q(N96) );
  AND2X1 U8 ( .IN1(bra_off0[28]), .IN2(n2), .Q(N95) );
  AND2X1 U9 ( .IN1(bra_off0[27]), .IN2(n2), .Q(N94) );
  AND2X1 U10 ( .IN1(bra_off0[26]), .IN2(n2), .Q(N93) );
  AND2X1 U11 ( .IN1(bra_off0[25]), .IN2(n2), .Q(N92) );
  AND2X1 U12 ( .IN1(bra_off0[24]), .IN2(n2), .Q(N91) );
  AND2X1 U13 ( .IN1(bra_off0[23]), .IN2(n2), .Q(N90) );
  AND2X1 U14 ( .IN1(cur_pc0[6]), .IN2(n2), .Q(N9) );
  AND2X1 U15 ( .IN1(bra_off0[22]), .IN2(n2), .Q(N89) );
  AND2X1 U16 ( .IN1(bra_off0[21]), .IN2(n2), .Q(N88) );
  AND2X1 U17 ( .IN1(bra_off0[20]), .IN2(n2), .Q(N87) );
  AND2X1 U18 ( .IN1(bra_off0[19]), .IN2(n2), .Q(N86) );
  AND2X1 U19 ( .IN1(bra_off0[18]), .IN2(n2), .Q(N85) );
  AND2X1 U20 ( .IN1(bra_off0[17]), .IN2(n2), .Q(N84) );
  AND2X1 U21 ( .IN1(bra_off0[16]), .IN2(n16), .Q(N83) );
  AND2X1 U22 ( .IN1(bra_off0[15]), .IN2(n16), .Q(N82) );
  AND2X1 U23 ( .IN1(bra_off0[14]), .IN2(n16), .Q(N81) );
  AND2X1 U24 ( .IN1(bra_off0[13]), .IN2(n16), .Q(N80) );
  AND2X1 U25 ( .IN1(cur_pc0[5]), .IN2(n16), .Q(N8) );
  AND2X1 U26 ( .IN1(bra_off0[12]), .IN2(n16), .Q(N79) );
  AND2X1 U27 ( .IN1(bra_off0[11]), .IN2(n16), .Q(N78) );
  AND2X1 U28 ( .IN1(bra_off0[10]), .IN2(n16), .Q(N77) );
  AND2X1 U29 ( .IN1(bra_off0[9]), .IN2(n16), .Q(N76) );
  AND2X1 U30 ( .IN1(bra_off0[8]), .IN2(n16), .Q(N75) );
  AND2X1 U31 ( .IN1(bra_off0[7]), .IN2(n16), .Q(N74) );
  AND2X1 U32 ( .IN1(bra_off0[6]), .IN2(n16), .Q(N73) );
  AND2X1 U33 ( .IN1(bra_off0[5]), .IN2(n15), .Q(N72) );
  AND2X1 U34 ( .IN1(bra_off0[4]), .IN2(n15), .Q(N71) );
  AND2X1 U35 ( .IN1(bra_off0[3]), .IN2(n15), .Q(N70) );
  AND2X1 U36 ( .IN1(cur_pc0[4]), .IN2(n15), .Q(N7) );
  AND2X1 U37 ( .IN1(bra_off0[2]), .IN2(n15), .Q(N69) );
  AND2X1 U38 ( .IN1(bra_off0[1]), .IN2(n15), .Q(N68) );
  AND2X1 U39 ( .IN1(bra_off0[0]), .IN2(n15), .Q(N67) );
  AND2X1 U40 ( .IN1(next_pc0[31]), .IN2(n15), .Q(N66) );
  AND2X1 U41 ( .IN1(next_pc0[30]), .IN2(n15), .Q(N65) );
  AND2X1 U42 ( .IN1(next_pc0[29]), .IN2(n15), .Q(N64) );
  AND2X1 U43 ( .IN1(next_pc0[28]), .IN2(n15), .Q(N63) );
  AND2X1 U44 ( .IN1(next_pc0[27]), .IN2(n15), .Q(N62) );
  AND2X1 U45 ( .IN1(next_pc0[26]), .IN2(n14), .Q(N61) );
  AND2X1 U46 ( .IN1(next_pc0[25]), .IN2(n14), .Q(N60) );
  AND2X1 U47 ( .IN1(cur_pc0[3]), .IN2(n14), .Q(N6) );
  AND2X1 U48 ( .IN1(next_pc0[24]), .IN2(n14), .Q(N59) );
  AND2X1 U49 ( .IN1(next_pc0[23]), .IN2(n14), .Q(N58) );
  AND2X1 U50 ( .IN1(next_pc0[22]), .IN2(n14), .Q(N57) );
  AND2X1 U51 ( .IN1(next_pc0[21]), .IN2(n14), .Q(N56) );
  AND2X1 U52 ( .IN1(next_pc0[20]), .IN2(n14), .Q(N55) );
  AND2X1 U53 ( .IN1(next_pc0[19]), .IN2(n14), .Q(N54) );
  AND2X1 U54 ( .IN1(next_pc0[18]), .IN2(n14), .Q(N53) );
  AND2X1 U55 ( .IN1(next_pc0[17]), .IN2(n14), .Q(N52) );
  AND2X1 U56 ( .IN1(next_pc0[16]), .IN2(n14), .Q(N51) );
  AND2X1 U57 ( .IN1(next_pc0[15]), .IN2(n13), .Q(N50) );
  AND2X1 U58 ( .IN1(cur_pc0[2]), .IN2(n13), .Q(N5) );
  AND2X1 U59 ( .IN1(next_pc0[14]), .IN2(n13), .Q(N49) );
  AND2X1 U60 ( .IN1(next_pc0[13]), .IN2(n13), .Q(N48) );
  AND2X1 U61 ( .IN1(next_pc0[12]), .IN2(n13), .Q(N47) );
  AND2X1 U62 ( .IN1(next_pc0[11]), .IN2(n13), .Q(N46) );
  AND2X1 U63 ( .IN1(next_pc0[10]), .IN2(n13), .Q(N45) );
  AND2X1 U64 ( .IN1(next_pc0[9]), .IN2(n13), .Q(N44) );
  AND2X1 U65 ( .IN1(next_pc0[8]), .IN2(n13), .Q(N43) );
  AND2X1 U66 ( .IN1(next_pc0[7]), .IN2(n13), .Q(N42) );
  AND2X1 U67 ( .IN1(next_pc0[6]), .IN2(n13), .Q(N41) );
  AND2X1 U68 ( .IN1(next_pc0[5]), .IN2(n13), .Q(N40) );
  AND2X1 U69 ( .IN1(cur_pc0[1]), .IN2(n12), .Q(N4) );
  AND2X1 U70 ( .IN1(next_pc0[4]), .IN2(n12), .Q(N39) );
  AND2X1 U71 ( .IN1(next_pc0[3]), .IN2(n12), .Q(N38) );
  AND2X1 U72 ( .IN1(next_pc0[2]), .IN2(n12), .Q(N37) );
  AND2X1 U73 ( .IN1(next_pc0[1]), .IN2(n12), .Q(N36) );
  AND2X1 U74 ( .IN1(next_pc0[0]), .IN2(n12), .Q(N35) );
  AND2X1 U75 ( .IN1(cur_pc0[31]), .IN2(n12), .Q(N34) );
  AND2X1 U76 ( .IN1(cur_pc0[30]), .IN2(n12), .Q(N33) );
  AND2X1 U77 ( .IN1(cur_pc0[29]), .IN2(n12), .Q(N32) );
  AND2X1 U78 ( .IN1(cur_pc0[28]), .IN2(n12), .Q(N31) );
  AND2X1 U79 ( .IN1(cur_pc0[27]), .IN2(n12), .Q(N30) );
  AND2X1 U80 ( .IN1(cur_pc0[0]), .IN2(n12), .Q(N3) );
  AND2X1 U81 ( .IN1(cur_pc0[26]), .IN2(n11), .Q(N29) );
  AND2X1 U82 ( .IN1(cur_pc0[25]), .IN2(n11), .Q(N28) );
  AND2X1 U83 ( .IN1(cur_pc0[24]), .IN2(n11), .Q(N27) );
  AND2X1 U84 ( .IN1(cur_pc0[23]), .IN2(n11), .Q(N26) );
  AND2X1 U85 ( .IN1(cur_pc0[22]), .IN2(n11), .Q(N25) );
  AND2X1 U86 ( .IN1(cur_pc0[21]), .IN2(n11), .Q(N24) );
  AND2X1 U87 ( .IN1(cur_pc0[20]), .IN2(n11), .Q(N23) );
  AND2X1 U88 ( .IN1(cur_pc0[19]), .IN2(n11), .Q(N22) );
  AND2X1 U89 ( .IN1(cur_pc0[18]), .IN2(n11), .Q(N21) );
  AND2X1 U90 ( .IN1(cur_pc0[17]), .IN2(n11), .Q(N20) );
  AND2X1 U91 ( .IN1(reg_addr0[4]), .IN2(n11), .Q(N199) );
  AND2X1 U92 ( .IN1(reg_addr0[3]), .IN2(n11), .Q(N198) );
  AND2X1 U93 ( .IN1(reg_addr0[2]), .IN2(n10), .Q(N197) );
  AND2X1 U94 ( .IN1(reg_addr0[1]), .IN2(n10), .Q(N196) );
  AND2X1 U95 ( .IN1(reg_addr0[0]), .IN2(n10), .Q(N195) );
  AND2X1 U96 ( .IN1(mem_data0[31]), .IN2(n10), .Q(N194) );
  AND2X1 U97 ( .IN1(mem_data0[30]), .IN2(n10), .Q(N193) );
  AND2X1 U98 ( .IN1(mem_data0[29]), .IN2(n10), .Q(N192) );
  AND2X1 U99 ( .IN1(mem_data0[28]), .IN2(n10), .Q(N191) );
  AND2X1 U100 ( .IN1(mem_data0[27]), .IN2(n10), .Q(N190) );
  AND2X1 U101 ( .IN1(cur_pc0[16]), .IN2(n10), .Q(N19) );
  AND2X1 U102 ( .IN1(mem_data0[26]), .IN2(n10), .Q(N189) );
  AND2X1 U103 ( .IN1(mem_data0[25]), .IN2(n10), .Q(N188) );
  AND2X1 U104 ( .IN1(mem_data0[24]), .IN2(n10), .Q(N187) );
  AND2X1 U105 ( .IN1(mem_data0[23]), .IN2(n9), .Q(N186) );
  AND2X1 U106 ( .IN1(mem_data0[22]), .IN2(n9), .Q(N185) );
  AND2X1 U107 ( .IN1(mem_data0[21]), .IN2(n9), .Q(N184) );
  AND2X1 U108 ( .IN1(mem_data0[20]), .IN2(n9), .Q(N183) );
  AND2X1 U109 ( .IN1(mem_data0[19]), .IN2(n9), .Q(N182) );
  AND2X1 U110 ( .IN1(mem_data0[18]), .IN2(n9), .Q(N181) );
  AND2X1 U111 ( .IN1(mem_data0[17]), .IN2(n9), .Q(N180) );
  AND2X1 U112 ( .IN1(cur_pc0[15]), .IN2(n9), .Q(N18) );
  AND2X1 U113 ( .IN1(mem_data0[16]), .IN2(n9), .Q(N179) );
  AND2X1 U114 ( .IN1(mem_data0[15]), .IN2(n9), .Q(N178) );
  AND2X1 U115 ( .IN1(mem_data0[14]), .IN2(n9), .Q(N177) );
  AND2X1 U116 ( .IN1(mem_data0[13]), .IN2(n9), .Q(N176) );
  AND2X1 U117 ( .IN1(mem_data0[12]), .IN2(n8), .Q(N175) );
  AND2X1 U118 ( .IN1(mem_data0[11]), .IN2(n8), .Q(N174) );
  AND2X1 U119 ( .IN1(mem_data0[10]), .IN2(n8), .Q(N173) );
  AND2X1 U120 ( .IN1(mem_data0[9]), .IN2(n8), .Q(N172) );
  AND2X1 U121 ( .IN1(mem_data0[8]), .IN2(n8), .Q(N171) );
  AND2X1 U122 ( .IN1(mem_data0[7]), .IN2(n8), .Q(N170) );
  AND2X1 U123 ( .IN1(cur_pc0[14]), .IN2(n8), .Q(N17) );
  AND2X1 U124 ( .IN1(mem_data0[6]), .IN2(n8), .Q(N169) );
  AND2X1 U125 ( .IN1(mem_data0[5]), .IN2(n8), .Q(N168) );
  AND2X1 U126 ( .IN1(mem_data0[4]), .IN2(n8), .Q(N167) );
  AND2X1 U127 ( .IN1(mem_data0[3]), .IN2(n8), .Q(N166) );
  AND2X1 U128 ( .IN1(mem_data0[2]), .IN2(n8), .Q(N165) );
  AND2X1 U129 ( .IN1(mem_data0[1]), .IN2(n7), .Q(N164) );
  AND2X1 U130 ( .IN1(mem_data0[0]), .IN2(n7), .Q(N163) );
  AND2X1 U131 ( .IN1(opB0[31]), .IN2(n7), .Q(N162) );
  AND2X1 U132 ( .IN1(opB0[30]), .IN2(n7), .Q(N161) );
  AND2X1 U133 ( .IN1(opB0[29]), .IN2(n7), .Q(N160) );
  AND2X1 U134 ( .IN1(cur_pc0[13]), .IN2(n7), .Q(N16) );
  AND2X1 U135 ( .IN1(opB0[28]), .IN2(n7), .Q(N159) );
  AND2X1 U136 ( .IN1(opB0[27]), .IN2(n7), .Q(N158) );
  AND2X1 U137 ( .IN1(opB0[26]), .IN2(n7), .Q(N157) );
  AND2X1 U138 ( .IN1(opB0[25]), .IN2(n7), .Q(N156) );
  AND2X1 U139 ( .IN1(opB0[24]), .IN2(n7), .Q(N155) );
  AND2X1 U140 ( .IN1(opB0[23]), .IN2(n7), .Q(N154) );
  AND2X1 U141 ( .IN1(opB0[22]), .IN2(n6), .Q(N153) );
  AND2X1 U142 ( .IN1(opB0[21]), .IN2(n6), .Q(N152) );
  AND2X1 U143 ( .IN1(opB0[20]), .IN2(n6), .Q(N151) );
  AND2X1 U144 ( .IN1(opB0[19]), .IN2(n6), .Q(N150) );
  AND2X1 U145 ( .IN1(cur_pc0[12]), .IN2(n6), .Q(N15) );
  AND2X1 U146 ( .IN1(opB0[18]), .IN2(n6), .Q(N149) );
  AND2X1 U147 ( .IN1(opB0[17]), .IN2(n6), .Q(N148) );
  AND2X1 U148 ( .IN1(opB0[16]), .IN2(n6), .Q(N147) );
  AND2X1 U149 ( .IN1(opB0[15]), .IN2(n6), .Q(N146) );
  AND2X1 U150 ( .IN1(opB0[14]), .IN2(n6), .Q(N145) );
  AND2X1 U151 ( .IN1(opB0[13]), .IN2(n6), .Q(N144) );
  AND2X1 U152 ( .IN1(opB0[12]), .IN2(n6), .Q(N143) );
  AND2X1 U153 ( .IN1(opB0[11]), .IN2(n5), .Q(N142) );
  AND2X1 U154 ( .IN1(opB0[10]), .IN2(n5), .Q(N141) );
  AND2X1 U155 ( .IN1(opB0[9]), .IN2(n5), .Q(N140) );
  AND2X1 U156 ( .IN1(cur_pc0[11]), .IN2(n5), .Q(N14) );
  AND2X1 U157 ( .IN1(opB0[8]), .IN2(n5), .Q(N139) );
  AND2X1 U158 ( .IN1(opB0[7]), .IN2(n5), .Q(N138) );
  AND2X1 U159 ( .IN1(opB0[6]), .IN2(n5), .Q(N137) );
  AND2X1 U160 ( .IN1(opB0[5]), .IN2(n5), .Q(N136) );
  AND2X1 U161 ( .IN1(opB0[4]), .IN2(n5), .Q(N135) );
  AND2X1 U162 ( .IN1(opB0[3]), .IN2(n5), .Q(N134) );
  AND2X1 U163 ( .IN1(opB0[2]), .IN2(n5), .Q(N133) );
  AND2X1 U164 ( .IN1(opB0[1]), .IN2(n5), .Q(N132) );
  AND2X1 U165 ( .IN1(opB0[0]), .IN2(n4), .Q(N131) );
  AND2X1 U166 ( .IN1(opA0[31]), .IN2(n4), .Q(N130) );
  AND2X1 U167 ( .IN1(cur_pc0[10]), .IN2(n4), .Q(N13) );
  AND2X1 U168 ( .IN1(opA0[30]), .IN2(n4), .Q(N129) );
  AND2X1 U169 ( .IN1(opA0[29]), .IN2(n4), .Q(N128) );
  AND2X1 U170 ( .IN1(opA0[28]), .IN2(n4), .Q(N127) );
  AND2X1 U171 ( .IN1(opA0[27]), .IN2(n4), .Q(N126) );
  AND2X1 U172 ( .IN1(opA0[26]), .IN2(n4), .Q(N125) );
  AND2X1 U173 ( .IN1(opA0[25]), .IN2(n4), .Q(N124) );
  AND2X1 U174 ( .IN1(opA0[24]), .IN2(n4), .Q(N123) );
  AND2X1 U175 ( .IN1(opA0[23]), .IN2(n4), .Q(N122) );
  AND2X1 U176 ( .IN1(opA0[22]), .IN2(n4), .Q(N121) );
  AND2X1 U177 ( .IN1(opA0[21]), .IN2(n3), .Q(N120) );
  AND2X1 U178 ( .IN1(cur_pc0[9]), .IN2(n3), .Q(N12) );
  AND2X1 U179 ( .IN1(opA0[20]), .IN2(n3), .Q(N119) );
  AND2X1 U180 ( .IN1(opA0[19]), .IN2(n3), .Q(N118) );
  AND2X1 U181 ( .IN1(opA0[18]), .IN2(n3), .Q(N117) );
  AND2X1 U182 ( .IN1(opA0[17]), .IN2(n3), .Q(N116) );
  AND2X1 U183 ( .IN1(opA0[16]), .IN2(n3), .Q(N115) );
  AND2X1 U184 ( .IN1(opA0[15]), .IN2(n3), .Q(N114) );
  AND2X1 U185 ( .IN1(opA0[14]), .IN2(n3), .Q(N113) );
  AND2X1 U186 ( .IN1(opA0[13]), .IN2(n3), .Q(N112) );
  AND2X1 U187 ( .IN1(opA0[12]), .IN2(n3), .Q(N111) );
  AND2X1 U188 ( .IN1(opA0[11]), .IN2(n3), .Q(N110) );
  AND2X1 U189 ( .IN1(cur_pc0[8]), .IN2(n1), .Q(N11) );
  AND2X1 U190 ( .IN1(opA0[10]), .IN2(n1), .Q(N109) );
  AND2X1 U191 ( .IN1(opA0[9]), .IN2(n1), .Q(N108) );
  AND2X1 U192 ( .IN1(opA0[8]), .IN2(n1), .Q(N107) );
  AND2X1 U193 ( .IN1(opA0[7]), .IN2(n1), .Q(N106) );
  AND2X1 U194 ( .IN1(opA0[6]), .IN2(n1), .Q(N105) );
  AND2X1 U195 ( .IN1(opA0[5]), .IN2(n1), .Q(N104) );
  AND2X1 U196 ( .IN1(opA0[4]), .IN2(n1), .Q(N103) );
  AND2X1 U197 ( .IN1(opA0[3]), .IN2(n1), .Q(N102) );
  AND2X1 U198 ( .IN1(opA0[2]), .IN2(n1), .Q(N101) );
  AND2X1 U199 ( .IN1(opA0[1]), .IN2(n1), .Q(N100) );
  AND2X1 U200 ( .IN1(cur_pc0[7]), .IN2(n1), .Q(N10) );
  AND3X1 U201 ( .IN1(en), .IN2(n18), .IN3(nrst), .Q(n2) );
  INVX0 U3 ( .INP(n2), .ZN(n17) );
  INVX0 U202 ( .INP(n17), .ZN(n13) );
  INVX0 U203 ( .INP(n17), .ZN(n14) );
  INVX0 U204 ( .INP(n17), .ZN(n15) );
  INVX0 U205 ( .INP(n17), .ZN(n16) );
  INVX0 U206 ( .INP(n17), .ZN(n7) );
  INVX0 U207 ( .INP(n17), .ZN(n8) );
  INVX0 U208 ( .INP(n17), .ZN(n9) );
  INVX0 U209 ( .INP(n17), .ZN(n12) );
  INVX0 U210 ( .INP(n17), .ZN(n10) );
  INVX0 U211 ( .INP(n17), .ZN(n11) );
  INVX0 U212 ( .INP(n17), .ZN(n1) );
  INVX0 U213 ( .INP(n17), .ZN(n3) );
  INVX0 U214 ( .INP(n17), .ZN(n4) );
  INVX0 U215 ( .INP(n17), .ZN(n5) );
  INVX0 U216 ( .INP(n17), .ZN(n6) );
  INVX0 U217 ( .INP(flush), .ZN(n18) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  FADDX1 U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FADDX1 U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FADDX1 U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FADDX1 U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FADDX1 U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FADDX1 U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FADDX1 U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FADDX1 U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_31 ( .IN1(A[31]), .IN2(n2), .IN3(carry[31]), .Q(DIFF[31]) );
  INVX0 U1 ( .INP(B[1]), .ZN(n32) );
  NAND2X1 U2 ( .IN1(B[0]), .IN2(n1), .QN(carry[1]) );
  INVX0 U3 ( .INP(B[2]), .ZN(n31) );
  INVX0 U4 ( .INP(B[3]), .ZN(n30) );
  INVX0 U5 ( .INP(B[4]), .ZN(n29) );
  INVX0 U6 ( .INP(B[5]), .ZN(n28) );
  INVX0 U7 ( .INP(B[6]), .ZN(n27) );
  INVX0 U8 ( .INP(B[7]), .ZN(n26) );
  INVX0 U9 ( .INP(B[8]), .ZN(n25) );
  INVX0 U10 ( .INP(B[9]), .ZN(n24) );
  INVX0 U11 ( .INP(B[10]), .ZN(n23) );
  INVX0 U12 ( .INP(B[11]), .ZN(n22) );
  INVX0 U13 ( .INP(B[12]), .ZN(n21) );
  INVX0 U14 ( .INP(B[13]), .ZN(n20) );
  INVX0 U15 ( .INP(B[14]), .ZN(n19) );
  INVX0 U16 ( .INP(B[15]), .ZN(n18) );
  INVX0 U17 ( .INP(B[16]), .ZN(n17) );
  INVX0 U18 ( .INP(B[17]), .ZN(n16) );
  INVX0 U19 ( .INP(B[18]), .ZN(n15) );
  INVX0 U20 ( .INP(B[19]), .ZN(n14) );
  INVX0 U21 ( .INP(B[20]), .ZN(n13) );
  INVX0 U22 ( .INP(B[21]), .ZN(n12) );
  INVX0 U23 ( .INP(B[22]), .ZN(n11) );
  INVX0 U24 ( .INP(B[23]), .ZN(n10) );
  INVX0 U25 ( .INP(B[24]), .ZN(n9) );
  INVX0 U26 ( .INP(B[25]), .ZN(n8) );
  INVX0 U27 ( .INP(B[26]), .ZN(n7) );
  INVX0 U28 ( .INP(B[27]), .ZN(n6) );
  INVX0 U29 ( .INP(B[28]), .ZN(n5) );
  INVX0 U30 ( .INP(B[29]), .ZN(n4) );
  INVX0 U31 ( .INP(B[30]), .ZN(n3) );
  INVX0 U32 ( .INP(A[0]), .ZN(n1) );
  INVX0 U33 ( .INP(B[0]), .ZN(n33) );
  INVX0 U34 ( .INP(B[31]), .ZN(n2) );
  XOR2X1 U35 ( .IN1(n1), .IN2(n33), .Q(DIFF[0]) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_31 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry[31]), .Q(SUM[31]) );
  AND2X1 U1 ( .IN1(B[0]), .IN2(A[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module alu ( opA, opB, res, alu_code, z );
  input [31:0] opA;
  input [31:0] opB;
  output [31:0] res;
  input [6:0] alu_code;
  output z;
  wire   N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n13, n14, n15, n16, n17, n18, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  NOR4X0 U18 ( .IN1(n19), .IN2(n20), .IN3(n21), .IN4(n22), .QN(z) );
  OR4X1 U19 ( .IN1(res[23]), .IN2(res[24]), .IN3(res[25]), .IN4(res[26]), .Q(
        n22) );
  OR4X1 U20 ( .IN1(res[27]), .IN2(res[28]), .IN3(res[29]), .IN4(res[2]), .Q(
        n21) );
  NAND4X0 U21 ( .IN1(n86), .IN2(n85), .IN3(n23), .IN4(n24), .QN(n20) );
  NOR4X0 U22 ( .IN1(res[4]), .IN2(res[3]), .IN3(res[31]), .IN4(res[30]), .QN(
        n24) );
  NOR3X0 U23 ( .IN1(res[7]), .IN2(res[9]), .IN3(res[8]), .QN(n23) );
  OR4X1 U24 ( .IN1(n25), .IN2(n26), .IN3(n27), .IN4(n28), .Q(n19) );
  OR4X1 U25 ( .IN1(res[16]), .IN2(res[17]), .IN3(res[18]), .IN4(res[19]), .Q(
        n28) );
  OR4X1 U26 ( .IN1(res[1]), .IN2(res[20]), .IN3(res[21]), .IN4(res[22]), .Q(
        n27) );
  OR4X1 U27 ( .IN1(n29), .IN2(res[0]), .IN3(res[10]), .IN4(res[11]), .Q(n26)
         );
  AND3X1 U28 ( .IN1(n30), .IN2(n31), .IN3(n32), .Q(n29) );
  OR4X1 U29 ( .IN1(res[12]), .IN2(res[13]), .IN3(res[14]), .IN4(res[15]), .Q(
        n25) );
  AO22X1 U30 ( .IN1(N40), .IN2(n88), .IN3(N72), .IN4(n87), .Q(res[9]) );
  AO22X1 U31 ( .IN1(N39), .IN2(n88), .IN3(N71), .IN4(n87), .Q(res[8]) );
  AO22X1 U32 ( .IN1(N38), .IN2(n88), .IN3(N70), .IN4(n87), .Q(res[7]) );
  AO22X1 U33 ( .IN1(N37), .IN2(n88), .IN3(N69), .IN4(n87), .Q(res[6]) );
  AO22X1 U34 ( .IN1(N36), .IN2(n88), .IN3(N68), .IN4(n87), .Q(res[5]) );
  AO22X1 U35 ( .IN1(N35), .IN2(n88), .IN3(N67), .IN4(n87), .Q(res[4]) );
  AO22X1 U36 ( .IN1(N34), .IN2(n88), .IN3(N66), .IN4(n87), .Q(res[3]) );
  AO22X1 U37 ( .IN1(N62), .IN2(n88), .IN3(N94), .IN4(n87), .Q(res[31]) );
  AO22X1 U38 ( .IN1(N61), .IN2(n88), .IN3(N93), .IN4(n87), .Q(res[30]) );
  AO22X1 U39 ( .IN1(N33), .IN2(n88), .IN3(N65), .IN4(n87), .Q(res[2]) );
  AO22X1 U40 ( .IN1(N60), .IN2(n88), .IN3(N92), .IN4(n87), .Q(res[29]) );
  AO22X1 U41 ( .IN1(N59), .IN2(n88), .IN3(N91), .IN4(n87), .Q(res[28]) );
  AO22X1 U42 ( .IN1(N58), .IN2(n88), .IN3(N90), .IN4(n87), .Q(res[27]) );
  AO22X1 U43 ( .IN1(N57), .IN2(n88), .IN3(N89), .IN4(n87), .Q(res[26]) );
  AO22X1 U44 ( .IN1(N56), .IN2(n88), .IN3(N88), .IN4(n87), .Q(res[25]) );
  AO22X1 U45 ( .IN1(N55), .IN2(n88), .IN3(N87), .IN4(n87), .Q(res[24]) );
  AO22X1 U46 ( .IN1(N54), .IN2(n88), .IN3(N86), .IN4(n87), .Q(res[23]) );
  AO22X1 U47 ( .IN1(N53), .IN2(n88), .IN3(N85), .IN4(n87), .Q(res[22]) );
  AO22X1 U48 ( .IN1(N52), .IN2(n88), .IN3(N84), .IN4(n87), .Q(res[21]) );
  AO22X1 U49 ( .IN1(N51), .IN2(n88), .IN3(N83), .IN4(n87), .Q(res[20]) );
  AO22X1 U50 ( .IN1(N32), .IN2(n88), .IN3(N64), .IN4(n87), .Q(res[1]) );
  AO22X1 U51 ( .IN1(N50), .IN2(n88), .IN3(N82), .IN4(n87), .Q(res[19]) );
  AO22X1 U52 ( .IN1(N49), .IN2(n88), .IN3(N81), .IN4(n87), .Q(res[18]) );
  AO22X1 U53 ( .IN1(N48), .IN2(n88), .IN3(N80), .IN4(n87), .Q(res[17]) );
  AO22X1 U54 ( .IN1(N47), .IN2(n88), .IN3(N79), .IN4(n87), .Q(res[16]) );
  AO22X1 U55 ( .IN1(N46), .IN2(n88), .IN3(N78), .IN4(n87), .Q(res[15]) );
  AO22X1 U56 ( .IN1(N45), .IN2(n88), .IN3(N77), .IN4(n87), .Q(res[14]) );
  AO22X1 U57 ( .IN1(N44), .IN2(n88), .IN3(N76), .IN4(n87), .Q(res[13]) );
  AO22X1 U58 ( .IN1(N43), .IN2(n88), .IN3(N75), .IN4(n87), .Q(res[12]) );
  AO22X1 U59 ( .IN1(N42), .IN2(n88), .IN3(N74), .IN4(n87), .Q(res[11]) );
  AO22X1 U60 ( .IN1(N41), .IN2(n88), .IN3(N73), .IN4(n87), .Q(res[10]) );
  AO222X1 U61 ( .IN1(N63), .IN2(n87), .IN3(n35), .IN4(N95), .IN5(N31), .IN6(
        n88), .Q(res[0]) );
  NAND4X0 U62 ( .IN1(alu_code[5]), .IN2(n34), .IN3(n90), .IN4(n89), .QN(n31)
         );
  AND2X1 U63 ( .IN1(n34), .IN2(n33), .Q(n35) );
  NAND4X0 U64 ( .IN1(alu_code[5]), .IN2(alu_code[1]), .IN3(n34), .IN4(n89), 
        .QN(n30) );
  NOR4X0 U65 ( .IN1(alu_code[2]), .IN2(alu_code[0]), .IN3(alu_code[6]), .IN4(
        alu_code[4]), .QN(n34) );
  alu_DW01_sub_0 sub_768 ( .A(opA), .B(opB), .CI(1'b0), .DIFF({N94, N93, N92, 
        N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, 
        N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63}) );
  alu_DW01_add_0 add_765 ( .A(opA), .B(opB), .CI(1'b0), .SUM({N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31}) );
  INVX0 U2 ( .INP(res[5]), .ZN(n86) );
  INVX0 U3 ( .INP(res[6]), .ZN(n85) );
  INVX0 U5 ( .INP(n30), .ZN(n87) );
  INVX0 U6 ( .INP(n31), .ZN(n88) );
  INVX0 U7 ( .INP(opA[3]), .ZN(n56) );
  INVX0 U8 ( .INP(opA[8]), .ZN(n61) );
  INVX0 U10 ( .INP(opA[14]), .ZN(n67) );
  INVX0 U11 ( .INP(opA[17]), .ZN(n70) );
  INVX0 U12 ( .INP(opA[20]), .ZN(n73) );
  INVX0 U13 ( .INP(opA[23]), .ZN(n76) );
  INVX0 U14 ( .INP(opA[26]), .ZN(n79) );
  INVX0 U15 ( .INP(opA[4]), .ZN(n57) );
  INVX0 U16 ( .INP(opA[1]), .ZN(n54) );
  NAND2X1 U17 ( .IN1(n33), .IN2(n34), .QN(n32) );
  INVX0 U66 ( .INP(opA[5]), .ZN(n58) );
  INVX0 U67 ( .INP(opA[11]), .ZN(n64) );
  INVX0 U68 ( .INP(opA[29]), .ZN(n82) );
  INVX0 U69 ( .INP(opB[31]), .ZN(n84) );
  INVX0 U70 ( .INP(opB[0]), .ZN(n53) );
  INVX0 U71 ( .INP(opA[2]), .ZN(n55) );
  INVX0 U72 ( .INP(opA[13]), .ZN(n66) );
  INVX0 U73 ( .INP(opA[15]), .ZN(n68) );
  INVX0 U74 ( .INP(opA[7]), .ZN(n60) );
  INVX0 U75 ( .INP(opA[19]), .ZN(n72) );
  INVX0 U76 ( .INP(opA[9]), .ZN(n62) );
  INVX0 U77 ( .INP(opA[10]), .ZN(n63) );
  INVX0 U78 ( .INP(opA[12]), .ZN(n65) );
  INVX0 U79 ( .INP(opA[16]), .ZN(n69) );
  INVX0 U80 ( .INP(opA[6]), .ZN(n59) );
  INVX0 U81 ( .INP(opA[18]), .ZN(n71) );
  NOR2X0 U82 ( .IN1(n89), .IN2(n90), .QN(n33) );
  INVX0 U83 ( .INP(opA[21]), .ZN(n74) );
  INVX0 U84 ( .INP(opA[25]), .ZN(n78) );
  INVX0 U85 ( .INP(opA[27]), .ZN(n80) );
  INVX0 U86 ( .INP(opA[22]), .ZN(n75) );
  INVX0 U87 ( .INP(opA[24]), .ZN(n77) );
  INVX0 U88 ( .INP(opA[28]), .ZN(n81) );
  INVX0 U89 ( .INP(opA[30]), .ZN(n83) );
  INVX0 U90 ( .INP(alu_code[1]), .ZN(n90) );
  INVX0 U91 ( .INP(alu_code[3]), .ZN(n89) );
  AND2X1 U92 ( .IN1(n83), .IN2(opB[30]), .Q(n51) );
  NOR2X0 U93 ( .IN1(n53), .IN2(opA[0]), .QN(n1) );
  AND2X1 U94 ( .IN1(n54), .IN2(n1), .Q(n2) );
  OA222X1 U95 ( .IN1(opB[2]), .IN2(n55), .IN3(opB[1]), .IN4(n2), .IN5(n1), 
        .IN6(n54), .Q(n3) );
  AO221X1 U96 ( .IN1(opB[2]), .IN2(n55), .IN3(opB[3]), .IN4(n56), .IN5(n3), 
        .Q(n4) );
  OA221X1 U97 ( .IN1(opB[4]), .IN2(n57), .IN3(opB[3]), .IN4(n56), .IN5(n4), 
        .Q(n5) );
  AO221X1 U98 ( .IN1(opB[4]), .IN2(n57), .IN3(opB[5]), .IN4(n58), .IN5(n5), 
        .Q(n6) );
  OA221X1 U99 ( .IN1(opB[6]), .IN2(n59), .IN3(opB[5]), .IN4(n58), .IN5(n6), 
        .Q(n7) );
  AO221X1 U100 ( .IN1(opB[6]), .IN2(n59), .IN3(opB[7]), .IN4(n60), .IN5(n7), 
        .Q(n8) );
  OA221X1 U101 ( .IN1(opB[8]), .IN2(n61), .IN3(opB[7]), .IN4(n60), .IN5(n8), 
        .Q(n9) );
  AO221X1 U102 ( .IN1(opB[8]), .IN2(n61), .IN3(opB[9]), .IN4(n62), .IN5(n9), 
        .Q(n10) );
  OA221X1 U103 ( .IN1(opB[9]), .IN2(n62), .IN3(opB[10]), .IN4(n63), .IN5(n10), 
        .Q(n13) );
  AO221X1 U104 ( .IN1(opB[10]), .IN2(n63), .IN3(opB[11]), .IN4(n64), .IN5(n13), 
        .Q(n14) );
  OA221X1 U105 ( .IN1(opB[12]), .IN2(n65), .IN3(opB[11]), .IN4(n64), .IN5(n14), 
        .Q(n15) );
  AO221X1 U106 ( .IN1(opB[12]), .IN2(n65), .IN3(opB[13]), .IN4(n66), .IN5(n15), 
        .Q(n16) );
  OA221X1 U107 ( .IN1(opB[14]), .IN2(n67), .IN3(opB[13]), .IN4(n66), .IN5(n16), 
        .Q(n17) );
  AO221X1 U108 ( .IN1(opB[14]), .IN2(n67), .IN3(opB[15]), .IN4(n68), .IN5(n17), 
        .Q(n18) );
  OA221X1 U109 ( .IN1(opB[16]), .IN2(n69), .IN3(opB[15]), .IN4(n68), .IN5(n18), 
        .Q(n36) );
  AO221X1 U110 ( .IN1(opB[16]), .IN2(n69), .IN3(opB[17]), .IN4(n70), .IN5(n36), 
        .Q(n37) );
  OA221X1 U111 ( .IN1(opB[18]), .IN2(n71), .IN3(opB[17]), .IN4(n70), .IN5(n37), 
        .Q(n38) );
  AO221X1 U112 ( .IN1(opB[18]), .IN2(n71), .IN3(opB[19]), .IN4(n72), .IN5(n38), 
        .Q(n39) );
  OA221X1 U113 ( .IN1(opB[20]), .IN2(n73), .IN3(opB[19]), .IN4(n72), .IN5(n39), 
        .Q(n40) );
  AO221X1 U114 ( .IN1(opB[20]), .IN2(n73), .IN3(opB[21]), .IN4(n74), .IN5(n40), 
        .Q(n41) );
  OA221X1 U115 ( .IN1(opB[22]), .IN2(n75), .IN3(opB[21]), .IN4(n74), .IN5(n41), 
        .Q(n42) );
  AO221X1 U116 ( .IN1(opB[22]), .IN2(n75), .IN3(opB[23]), .IN4(n76), .IN5(n42), 
        .Q(n43) );
  OA221X1 U117 ( .IN1(opB[24]), .IN2(n77), .IN3(opB[23]), .IN4(n76), .IN5(n43), 
        .Q(n44) );
  AO221X1 U118 ( .IN1(opB[24]), .IN2(n77), .IN3(opB[25]), .IN4(n78), .IN5(n44), 
        .Q(n45) );
  OA221X1 U119 ( .IN1(opB[26]), .IN2(n79), .IN3(opB[25]), .IN4(n78), .IN5(n45), 
        .Q(n46) );
  AO221X1 U120 ( .IN1(opB[26]), .IN2(n79), .IN3(opB[27]), .IN4(n80), .IN5(n46), 
        .Q(n47) );
  OA221X1 U121 ( .IN1(opB[28]), .IN2(n81), .IN3(opB[27]), .IN4(n80), .IN5(n47), 
        .Q(n48) );
  AO221X1 U122 ( .IN1(opB[28]), .IN2(n81), .IN3(opB[29]), .IN4(n82), .IN5(n48), 
        .Q(n49) );
  OA221X1 U123 ( .IN1(opB[30]), .IN2(n83), .IN3(opB[29]), .IN4(n82), .IN5(n49), 
        .Q(n50) );
  OA22X1 U124 ( .IN1(opA[31]), .IN2(n84), .IN3(n51), .IN4(n50), .Q(n52) );
  AO21X1 U125 ( .IN1(opA[31]), .IN2(n84), .IN3(n52), .Q(N95) );
endmodule


module exe_mem_reg ( clk, nrst, cur_pc0, next_pc0, alu_out0, mem_data0, 
        reg_addr0, cur_pc, next_pc, alu_out, mem_data, reg_addr );
  input [31:0] cur_pc0;
  input [31:0] next_pc0;
  input [31:0] alu_out0;
  input [31:0] mem_data0;
  input [4:0] reg_addr0;
  output [31:0] cur_pc;
  output [31:0] next_pc;
  output [31:0] alu_out;
  output [31:0] mem_data;
  output [4:0] reg_addr;
  input clk, nrst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  DFFX1 \mem_data_reg[31]  ( .D(N130), .CLK(clk), .Q(mem_data[31]) );
  DFFX1 \mem_data_reg[30]  ( .D(N129), .CLK(clk), .Q(mem_data[30]) );
  DFFX1 \mem_data_reg[29]  ( .D(N128), .CLK(clk), .Q(mem_data[29]) );
  DFFX1 \mem_data_reg[28]  ( .D(N127), .CLK(clk), .Q(mem_data[28]) );
  DFFX1 \mem_data_reg[27]  ( .D(N126), .CLK(clk), .Q(mem_data[27]) );
  DFFX1 \mem_data_reg[26]  ( .D(N125), .CLK(clk), .Q(mem_data[26]) );
  DFFX1 \mem_data_reg[25]  ( .D(N124), .CLK(clk), .Q(mem_data[25]) );
  DFFX1 \mem_data_reg[24]  ( .D(N123), .CLK(clk), .Q(mem_data[24]) );
  DFFX1 \mem_data_reg[23]  ( .D(N122), .CLK(clk), .Q(mem_data[23]) );
  DFFX1 \mem_data_reg[22]  ( .D(N121), .CLK(clk), .Q(mem_data[22]) );
  DFFX1 \mem_data_reg[21]  ( .D(N120), .CLK(clk), .Q(mem_data[21]) );
  DFFX1 \mem_data_reg[20]  ( .D(N119), .CLK(clk), .Q(mem_data[20]) );
  DFFX1 \mem_data_reg[19]  ( .D(N118), .CLK(clk), .Q(mem_data[19]) );
  DFFX1 \mem_data_reg[18]  ( .D(N117), .CLK(clk), .Q(mem_data[18]) );
  DFFX1 \mem_data_reg[17]  ( .D(N116), .CLK(clk), .Q(mem_data[17]) );
  DFFX1 \mem_data_reg[16]  ( .D(N115), .CLK(clk), .Q(mem_data[16]) );
  DFFX1 \mem_data_reg[15]  ( .D(N114), .CLK(clk), .Q(mem_data[15]) );
  DFFX1 \mem_data_reg[14]  ( .D(N113), .CLK(clk), .Q(mem_data[14]) );
  DFFX1 \mem_data_reg[13]  ( .D(N112), .CLK(clk), .Q(mem_data[13]) );
  DFFX1 \mem_data_reg[12]  ( .D(N111), .CLK(clk), .Q(mem_data[12]) );
  DFFX1 \mem_data_reg[11]  ( .D(N110), .CLK(clk), .Q(mem_data[11]) );
  DFFX1 \mem_data_reg[10]  ( .D(N109), .CLK(clk), .Q(mem_data[10]) );
  DFFX1 \mem_data_reg[9]  ( .D(N108), .CLK(clk), .Q(mem_data[9]) );
  DFFX1 \mem_data_reg[8]  ( .D(N107), .CLK(clk), .Q(mem_data[8]) );
  DFFX1 \mem_data_reg[7]  ( .D(N106), .CLK(clk), .Q(mem_data[7]) );
  DFFX1 \mem_data_reg[6]  ( .D(N105), .CLK(clk), .Q(mem_data[6]) );
  DFFX1 \mem_data_reg[5]  ( .D(N104), .CLK(clk), .Q(mem_data[5]) );
  DFFX1 \mem_data_reg[4]  ( .D(N103), .CLK(clk), .Q(mem_data[4]) );
  DFFX1 \mem_data_reg[3]  ( .D(N102), .CLK(clk), .Q(mem_data[3]) );
  DFFX1 \mem_data_reg[2]  ( .D(N101), .CLK(clk), .Q(mem_data[2]) );
  DFFX1 \mem_data_reg[1]  ( .D(N100), .CLK(clk), .Q(mem_data[1]) );
  DFFX1 \mem_data_reg[0]  ( .D(N99), .CLK(clk), .Q(mem_data[0]) );
  DFFX1 \reg_addr_reg[4]  ( .D(N135), .CLK(clk), .Q(reg_addr[4]) );
  DFFX1 \reg_addr_reg[3]  ( .D(N134), .CLK(clk), .Q(reg_addr[3]) );
  DFFX1 \reg_addr_reg[2]  ( .D(N133), .CLK(clk), .Q(reg_addr[2]) );
  DFFX1 \reg_addr_reg[1]  ( .D(N132), .CLK(clk), .Q(reg_addr[1]) );
  DFFX1 \reg_addr_reg[0]  ( .D(N131), .CLK(clk), .Q(reg_addr[0]) );
  DFFX1 \cur_pc_reg[31]  ( .D(N34), .CLK(clk), .Q(cur_pc[31]) );
  DFFX1 \cur_pc_reg[30]  ( .D(N33), .CLK(clk), .Q(cur_pc[30]) );
  DFFX1 \cur_pc_reg[29]  ( .D(N32), .CLK(clk), .Q(cur_pc[29]) );
  DFFX1 \cur_pc_reg[28]  ( .D(N31), .CLK(clk), .Q(cur_pc[28]) );
  DFFX1 \cur_pc_reg[27]  ( .D(N30), .CLK(clk), .Q(cur_pc[27]) );
  DFFX1 \cur_pc_reg[26]  ( .D(N29), .CLK(clk), .Q(cur_pc[26]) );
  DFFX1 \cur_pc_reg[25]  ( .D(N28), .CLK(clk), .Q(cur_pc[25]) );
  DFFX1 \cur_pc_reg[24]  ( .D(N27), .CLK(clk), .Q(cur_pc[24]) );
  DFFX1 \cur_pc_reg[23]  ( .D(N26), .CLK(clk), .Q(cur_pc[23]) );
  DFFX1 \cur_pc_reg[22]  ( .D(N25), .CLK(clk), .Q(cur_pc[22]) );
  DFFX1 \cur_pc_reg[21]  ( .D(N24), .CLK(clk), .Q(cur_pc[21]) );
  DFFX1 \cur_pc_reg[20]  ( .D(N23), .CLK(clk), .Q(cur_pc[20]) );
  DFFX1 \cur_pc_reg[19]  ( .D(N22), .CLK(clk), .Q(cur_pc[19]) );
  DFFX1 \cur_pc_reg[18]  ( .D(N21), .CLK(clk), .Q(cur_pc[18]) );
  DFFX1 \cur_pc_reg[17]  ( .D(N20), .CLK(clk), .Q(cur_pc[17]) );
  DFFX1 \cur_pc_reg[16]  ( .D(N19), .CLK(clk), .Q(cur_pc[16]) );
  DFFX1 \cur_pc_reg[15]  ( .D(N18), .CLK(clk), .Q(cur_pc[15]) );
  DFFX1 \cur_pc_reg[14]  ( .D(N17), .CLK(clk), .Q(cur_pc[14]) );
  DFFX1 \cur_pc_reg[13]  ( .D(N16), .CLK(clk), .Q(cur_pc[13]) );
  DFFX1 \cur_pc_reg[12]  ( .D(N15), .CLK(clk), .Q(cur_pc[12]) );
  DFFX1 \cur_pc_reg[11]  ( .D(N14), .CLK(clk), .Q(cur_pc[11]) );
  DFFX1 \cur_pc_reg[10]  ( .D(N13), .CLK(clk), .Q(cur_pc[10]) );
  DFFX1 \cur_pc_reg[9]  ( .D(N12), .CLK(clk), .Q(cur_pc[9]) );
  DFFX1 \cur_pc_reg[8]  ( .D(N11), .CLK(clk), .Q(cur_pc[8]) );
  DFFX1 \cur_pc_reg[7]  ( .D(N10), .CLK(clk), .Q(cur_pc[7]) );
  DFFX1 \cur_pc_reg[6]  ( .D(N9), .CLK(clk), .Q(cur_pc[6]) );
  DFFX1 \cur_pc_reg[5]  ( .D(N8), .CLK(clk), .Q(cur_pc[5]) );
  DFFX1 \cur_pc_reg[4]  ( .D(N7), .CLK(clk), .Q(cur_pc[4]) );
  DFFX1 \cur_pc_reg[3]  ( .D(N6), .CLK(clk), .Q(cur_pc[3]) );
  DFFX1 \cur_pc_reg[2]  ( .D(N5), .CLK(clk), .Q(cur_pc[2]) );
  DFFX1 \cur_pc_reg[1]  ( .D(N4), .CLK(clk), .Q(cur_pc[1]) );
  DFFX1 \cur_pc_reg[0]  ( .D(N3), .CLK(clk), .Q(cur_pc[0]) );
  DFFX1 \next_pc_reg[31]  ( .D(N66), .CLK(clk), .Q(next_pc[31]) );
  DFFX1 \next_pc_reg[30]  ( .D(N65), .CLK(clk), .Q(next_pc[30]) );
  DFFX1 \next_pc_reg[29]  ( .D(N64), .CLK(clk), .Q(next_pc[29]) );
  DFFX1 \next_pc_reg[28]  ( .D(N63), .CLK(clk), .Q(next_pc[28]) );
  DFFX1 \next_pc_reg[27]  ( .D(N62), .CLK(clk), .Q(next_pc[27]) );
  DFFX1 \next_pc_reg[26]  ( .D(N61), .CLK(clk), .Q(next_pc[26]) );
  DFFX1 \next_pc_reg[25]  ( .D(N60), .CLK(clk), .Q(next_pc[25]) );
  DFFX1 \next_pc_reg[24]  ( .D(N59), .CLK(clk), .Q(next_pc[24]) );
  DFFX1 \next_pc_reg[23]  ( .D(N58), .CLK(clk), .Q(next_pc[23]) );
  DFFX1 \next_pc_reg[22]  ( .D(N57), .CLK(clk), .Q(next_pc[22]) );
  DFFX1 \next_pc_reg[21]  ( .D(N56), .CLK(clk), .Q(next_pc[21]) );
  DFFX1 \next_pc_reg[20]  ( .D(N55), .CLK(clk), .Q(next_pc[20]) );
  DFFX1 \next_pc_reg[19]  ( .D(N54), .CLK(clk), .Q(next_pc[19]) );
  DFFX1 \next_pc_reg[18]  ( .D(N53), .CLK(clk), .Q(next_pc[18]) );
  DFFX1 \next_pc_reg[17]  ( .D(N52), .CLK(clk), .Q(next_pc[17]) );
  DFFX1 \next_pc_reg[16]  ( .D(N51), .CLK(clk), .Q(next_pc[16]) );
  DFFX1 \next_pc_reg[15]  ( .D(N50), .CLK(clk), .Q(next_pc[15]) );
  DFFX1 \next_pc_reg[14]  ( .D(N49), .CLK(clk), .Q(next_pc[14]) );
  DFFX1 \next_pc_reg[13]  ( .D(N48), .CLK(clk), .Q(next_pc[13]) );
  DFFX1 \next_pc_reg[12]  ( .D(N47), .CLK(clk), .Q(next_pc[12]) );
  DFFX1 \next_pc_reg[11]  ( .D(N46), .CLK(clk), .Q(next_pc[11]) );
  DFFX1 \next_pc_reg[10]  ( .D(N45), .CLK(clk), .Q(next_pc[10]) );
  DFFX1 \next_pc_reg[9]  ( .D(N44), .CLK(clk), .Q(next_pc[9]) );
  DFFX1 \next_pc_reg[8]  ( .D(N43), .CLK(clk), .Q(next_pc[8]) );
  DFFX1 \next_pc_reg[7]  ( .D(N42), .CLK(clk), .Q(next_pc[7]) );
  DFFX1 \next_pc_reg[6]  ( .D(N41), .CLK(clk), .Q(next_pc[6]) );
  DFFX1 \next_pc_reg[5]  ( .D(N40), .CLK(clk), .Q(next_pc[5]) );
  DFFX1 \next_pc_reg[4]  ( .D(N39), .CLK(clk), .Q(next_pc[4]) );
  DFFX1 \next_pc_reg[3]  ( .D(N38), .CLK(clk), .Q(next_pc[3]) );
  DFFX1 \next_pc_reg[2]  ( .D(N37), .CLK(clk), .Q(next_pc[2]) );
  DFFX1 \next_pc_reg[1]  ( .D(N36), .CLK(clk), .Q(next_pc[1]) );
  DFFX1 \next_pc_reg[0]  ( .D(N35), .CLK(clk), .Q(next_pc[0]) );
  DFFX1 \alu_out_reg[31]  ( .D(N98), .CLK(clk), .Q(alu_out[31]) );
  DFFX1 \alu_out_reg[30]  ( .D(N97), .CLK(clk), .Q(alu_out[30]) );
  DFFX1 \alu_out_reg[29]  ( .D(N96), .CLK(clk), .Q(alu_out[29]) );
  DFFX1 \alu_out_reg[28]  ( .D(N95), .CLK(clk), .Q(alu_out[28]) );
  DFFX1 \alu_out_reg[27]  ( .D(N94), .CLK(clk), .Q(alu_out[27]) );
  DFFX1 \alu_out_reg[26]  ( .D(N93), .CLK(clk), .Q(alu_out[26]) );
  DFFX1 \alu_out_reg[25]  ( .D(N92), .CLK(clk), .Q(alu_out[25]) );
  DFFX1 \alu_out_reg[24]  ( .D(N91), .CLK(clk), .Q(alu_out[24]) );
  DFFX1 \alu_out_reg[23]  ( .D(N90), .CLK(clk), .Q(alu_out[23]) );
  DFFX1 \alu_out_reg[22]  ( .D(N89), .CLK(clk), .Q(alu_out[22]) );
  DFFX1 \alu_out_reg[21]  ( .D(N88), .CLK(clk), .Q(alu_out[21]) );
  DFFX1 \alu_out_reg[20]  ( .D(N87), .CLK(clk), .Q(alu_out[20]) );
  DFFX1 \alu_out_reg[19]  ( .D(N86), .CLK(clk), .Q(alu_out[19]) );
  DFFX1 \alu_out_reg[18]  ( .D(N85), .CLK(clk), .Q(alu_out[18]) );
  DFFX1 \alu_out_reg[17]  ( .D(N84), .CLK(clk), .Q(alu_out[17]) );
  DFFX1 \alu_out_reg[16]  ( .D(N83), .CLK(clk), .Q(alu_out[16]) );
  DFFX1 \alu_out_reg[15]  ( .D(N82), .CLK(clk), .Q(alu_out[15]) );
  DFFX1 \alu_out_reg[14]  ( .D(N81), .CLK(clk), .Q(alu_out[14]) );
  DFFX1 \alu_out_reg[13]  ( .D(N80), .CLK(clk), .Q(alu_out[13]) );
  DFFX1 \alu_out_reg[12]  ( .D(N79), .CLK(clk), .Q(alu_out[12]) );
  DFFX1 \alu_out_reg[11]  ( .D(N78), .CLK(clk), .Q(alu_out[11]) );
  DFFX1 \alu_out_reg[10]  ( .D(N77), .CLK(clk), .Q(alu_out[10]) );
  DFFX1 \alu_out_reg[9]  ( .D(N76), .CLK(clk), .Q(alu_out[9]) );
  DFFX1 \alu_out_reg[8]  ( .D(N75), .CLK(clk), .Q(alu_out[8]) );
  DFFX1 \alu_out_reg[7]  ( .D(N74), .CLK(clk), .Q(alu_out[7]) );
  DFFX1 \alu_out_reg[6]  ( .D(N73), .CLK(clk), .Q(alu_out[6]) );
  DFFX1 \alu_out_reg[5]  ( .D(N72), .CLK(clk), .Q(alu_out[5]) );
  DFFX1 \alu_out_reg[4]  ( .D(N71), .CLK(clk), .Q(alu_out[4]) );
  DFFX1 \alu_out_reg[3]  ( .D(N70), .CLK(clk), .Q(alu_out[3]) );
  DFFX1 \alu_out_reg[2]  ( .D(N69), .CLK(clk), .Q(alu_out[2]) );
  DFFX1 \alu_out_reg[1]  ( .D(N68), .CLK(clk), .Q(alu_out[1]) );
  DFFX1 \alu_out_reg[0]  ( .D(N67), .CLK(clk), .Q(alu_out[0]) );
  AND2X1 U3 ( .IN1(nrst), .IN2(mem_data0[0]), .Q(N99) );
  AND2X1 U4 ( .IN1(alu_out0[31]), .IN2(n11), .Q(N98) );
  AND2X1 U5 ( .IN1(alu_out0[30]), .IN2(n11), .Q(N97) );
  AND2X1 U6 ( .IN1(alu_out0[29]), .IN2(n11), .Q(N96) );
  AND2X1 U7 ( .IN1(alu_out0[28]), .IN2(n11), .Q(N95) );
  AND2X1 U8 ( .IN1(alu_out0[27]), .IN2(n11), .Q(N94) );
  AND2X1 U9 ( .IN1(alu_out0[26]), .IN2(n11), .Q(N93) );
  AND2X1 U10 ( .IN1(alu_out0[25]), .IN2(n11), .Q(N92) );
  AND2X1 U11 ( .IN1(alu_out0[24]), .IN2(n11), .Q(N91) );
  AND2X1 U12 ( .IN1(alu_out0[23]), .IN2(n11), .Q(N90) );
  AND2X1 U13 ( .IN1(cur_pc0[6]), .IN2(n11), .Q(N9) );
  AND2X1 U14 ( .IN1(alu_out0[22]), .IN2(n11), .Q(N89) );
  AND2X1 U15 ( .IN1(alu_out0[21]), .IN2(n11), .Q(N88) );
  AND2X1 U16 ( .IN1(alu_out0[20]), .IN2(n10), .Q(N87) );
  AND2X1 U17 ( .IN1(alu_out0[19]), .IN2(n10), .Q(N86) );
  AND2X1 U18 ( .IN1(alu_out0[18]), .IN2(n10), .Q(N85) );
  AND2X1 U19 ( .IN1(alu_out0[17]), .IN2(n10), .Q(N84) );
  AND2X1 U20 ( .IN1(alu_out0[16]), .IN2(n10), .Q(N83) );
  AND2X1 U21 ( .IN1(alu_out0[15]), .IN2(n10), .Q(N82) );
  AND2X1 U22 ( .IN1(alu_out0[14]), .IN2(n10), .Q(N81) );
  AND2X1 U23 ( .IN1(alu_out0[13]), .IN2(n10), .Q(N80) );
  AND2X1 U24 ( .IN1(cur_pc0[5]), .IN2(n10), .Q(N8) );
  AND2X1 U25 ( .IN1(alu_out0[12]), .IN2(n10), .Q(N79) );
  AND2X1 U26 ( .IN1(alu_out0[11]), .IN2(n10), .Q(N78) );
  AND2X1 U27 ( .IN1(alu_out0[10]), .IN2(n10), .Q(N77) );
  AND2X1 U28 ( .IN1(alu_out0[9]), .IN2(n9), .Q(N76) );
  AND2X1 U29 ( .IN1(alu_out0[8]), .IN2(n9), .Q(N75) );
  AND2X1 U30 ( .IN1(alu_out0[7]), .IN2(n9), .Q(N74) );
  AND2X1 U31 ( .IN1(alu_out0[6]), .IN2(n9), .Q(N73) );
  AND2X1 U32 ( .IN1(alu_out0[5]), .IN2(n9), .Q(N72) );
  AND2X1 U33 ( .IN1(alu_out0[4]), .IN2(n9), .Q(N71) );
  AND2X1 U34 ( .IN1(alu_out0[3]), .IN2(n9), .Q(N70) );
  AND2X1 U35 ( .IN1(cur_pc0[4]), .IN2(n9), .Q(N7) );
  AND2X1 U36 ( .IN1(alu_out0[2]), .IN2(n9), .Q(N69) );
  AND2X1 U37 ( .IN1(alu_out0[1]), .IN2(n9), .Q(N68) );
  AND2X1 U38 ( .IN1(alu_out0[0]), .IN2(n9), .Q(N67) );
  AND2X1 U39 ( .IN1(next_pc0[31]), .IN2(n9), .Q(N66) );
  AND2X1 U40 ( .IN1(next_pc0[30]), .IN2(n8), .Q(N65) );
  AND2X1 U41 ( .IN1(next_pc0[29]), .IN2(n8), .Q(N64) );
  AND2X1 U42 ( .IN1(next_pc0[28]), .IN2(n8), .Q(N63) );
  AND2X1 U43 ( .IN1(next_pc0[27]), .IN2(n8), .Q(N62) );
  AND2X1 U44 ( .IN1(next_pc0[26]), .IN2(n8), .Q(N61) );
  AND2X1 U45 ( .IN1(next_pc0[25]), .IN2(n8), .Q(N60) );
  AND2X1 U46 ( .IN1(cur_pc0[3]), .IN2(n8), .Q(N6) );
  AND2X1 U47 ( .IN1(next_pc0[24]), .IN2(n8), .Q(N59) );
  AND2X1 U48 ( .IN1(next_pc0[23]), .IN2(n8), .Q(N58) );
  AND2X1 U49 ( .IN1(next_pc0[22]), .IN2(n8), .Q(N57) );
  AND2X1 U50 ( .IN1(next_pc0[21]), .IN2(n8), .Q(N56) );
  AND2X1 U51 ( .IN1(next_pc0[20]), .IN2(n8), .Q(N55) );
  AND2X1 U52 ( .IN1(next_pc0[19]), .IN2(n7), .Q(N54) );
  AND2X1 U53 ( .IN1(next_pc0[18]), .IN2(n7), .Q(N53) );
  AND2X1 U54 ( .IN1(next_pc0[17]), .IN2(n7), .Q(N52) );
  AND2X1 U55 ( .IN1(next_pc0[16]), .IN2(n7), .Q(N51) );
  AND2X1 U56 ( .IN1(next_pc0[15]), .IN2(n7), .Q(N50) );
  AND2X1 U57 ( .IN1(cur_pc0[2]), .IN2(n7), .Q(N5) );
  AND2X1 U58 ( .IN1(next_pc0[14]), .IN2(n7), .Q(N49) );
  AND2X1 U59 ( .IN1(next_pc0[13]), .IN2(n7), .Q(N48) );
  AND2X1 U60 ( .IN1(next_pc0[12]), .IN2(n7), .Q(N47) );
  AND2X1 U61 ( .IN1(next_pc0[11]), .IN2(n7), .Q(N46) );
  AND2X1 U62 ( .IN1(next_pc0[10]), .IN2(n7), .Q(N45) );
  AND2X1 U63 ( .IN1(next_pc0[9]), .IN2(n7), .Q(N44) );
  AND2X1 U64 ( .IN1(next_pc0[8]), .IN2(n6), .Q(N43) );
  AND2X1 U65 ( .IN1(next_pc0[7]), .IN2(n6), .Q(N42) );
  AND2X1 U66 ( .IN1(next_pc0[6]), .IN2(n6), .Q(N41) );
  AND2X1 U67 ( .IN1(next_pc0[5]), .IN2(n6), .Q(N40) );
  AND2X1 U68 ( .IN1(cur_pc0[1]), .IN2(n6), .Q(N4) );
  AND2X1 U69 ( .IN1(next_pc0[4]), .IN2(n6), .Q(N39) );
  AND2X1 U70 ( .IN1(next_pc0[3]), .IN2(n6), .Q(N38) );
  AND2X1 U71 ( .IN1(next_pc0[2]), .IN2(n6), .Q(N37) );
  AND2X1 U72 ( .IN1(next_pc0[1]), .IN2(n6), .Q(N36) );
  AND2X1 U73 ( .IN1(next_pc0[0]), .IN2(n6), .Q(N35) );
  AND2X1 U74 ( .IN1(cur_pc0[31]), .IN2(n6), .Q(N34) );
  AND2X1 U75 ( .IN1(cur_pc0[30]), .IN2(n6), .Q(N33) );
  AND2X1 U76 ( .IN1(cur_pc0[29]), .IN2(n5), .Q(N32) );
  AND2X1 U77 ( .IN1(cur_pc0[28]), .IN2(n5), .Q(N31) );
  AND2X1 U78 ( .IN1(cur_pc0[27]), .IN2(n5), .Q(N30) );
  AND2X1 U79 ( .IN1(cur_pc0[0]), .IN2(n5), .Q(N3) );
  AND2X1 U80 ( .IN1(cur_pc0[26]), .IN2(n5), .Q(N29) );
  AND2X1 U81 ( .IN1(cur_pc0[25]), .IN2(n5), .Q(N28) );
  AND2X1 U82 ( .IN1(cur_pc0[24]), .IN2(n5), .Q(N27) );
  AND2X1 U83 ( .IN1(cur_pc0[23]), .IN2(n5), .Q(N26) );
  AND2X1 U84 ( .IN1(cur_pc0[22]), .IN2(n5), .Q(N25) );
  AND2X1 U85 ( .IN1(cur_pc0[21]), .IN2(n5), .Q(N24) );
  AND2X1 U86 ( .IN1(cur_pc0[20]), .IN2(n5), .Q(N23) );
  AND2X1 U87 ( .IN1(cur_pc0[19]), .IN2(n5), .Q(N22) );
  AND2X1 U88 ( .IN1(cur_pc0[18]), .IN2(n4), .Q(N21) );
  AND2X1 U89 ( .IN1(cur_pc0[17]), .IN2(n4), .Q(N20) );
  AND2X1 U90 ( .IN1(cur_pc0[16]), .IN2(n4), .Q(N19) );
  AND2X1 U91 ( .IN1(cur_pc0[15]), .IN2(n4), .Q(N18) );
  AND2X1 U92 ( .IN1(cur_pc0[14]), .IN2(n4), .Q(N17) );
  AND2X1 U93 ( .IN1(cur_pc0[13]), .IN2(n4), .Q(N16) );
  AND2X1 U94 ( .IN1(cur_pc0[12]), .IN2(n4), .Q(N15) );
  AND2X1 U95 ( .IN1(cur_pc0[11]), .IN2(n4), .Q(N14) );
  AND2X1 U96 ( .IN1(reg_addr0[4]), .IN2(n4), .Q(N135) );
  AND2X1 U97 ( .IN1(reg_addr0[3]), .IN2(n4), .Q(N134) );
  AND2X1 U98 ( .IN1(reg_addr0[2]), .IN2(n4), .Q(N133) );
  AND2X1 U99 ( .IN1(reg_addr0[1]), .IN2(n4), .Q(N132) );
  AND2X1 U100 ( .IN1(reg_addr0[0]), .IN2(n3), .Q(N131) );
  AND2X1 U101 ( .IN1(mem_data0[31]), .IN2(n3), .Q(N130) );
  AND2X1 U102 ( .IN1(cur_pc0[10]), .IN2(n3), .Q(N13) );
  AND2X1 U103 ( .IN1(mem_data0[30]), .IN2(n3), .Q(N129) );
  AND2X1 U104 ( .IN1(mem_data0[29]), .IN2(n3), .Q(N128) );
  AND2X1 U105 ( .IN1(mem_data0[28]), .IN2(n3), .Q(N127) );
  AND2X1 U106 ( .IN1(mem_data0[27]), .IN2(n3), .Q(N126) );
  AND2X1 U107 ( .IN1(mem_data0[26]), .IN2(n3), .Q(N125) );
  AND2X1 U108 ( .IN1(mem_data0[25]), .IN2(n3), .Q(N124) );
  AND2X1 U109 ( .IN1(mem_data0[24]), .IN2(n3), .Q(N123) );
  AND2X1 U110 ( .IN1(mem_data0[23]), .IN2(n3), .Q(N122) );
  AND2X1 U111 ( .IN1(mem_data0[22]), .IN2(n3), .Q(N121) );
  AND2X1 U112 ( .IN1(mem_data0[21]), .IN2(n2), .Q(N120) );
  AND2X1 U113 ( .IN1(cur_pc0[9]), .IN2(n2), .Q(N12) );
  AND2X1 U114 ( .IN1(mem_data0[20]), .IN2(n2), .Q(N119) );
  AND2X1 U115 ( .IN1(mem_data0[19]), .IN2(n2), .Q(N118) );
  AND2X1 U116 ( .IN1(mem_data0[18]), .IN2(n2), .Q(N117) );
  AND2X1 U117 ( .IN1(mem_data0[17]), .IN2(n2), .Q(N116) );
  AND2X1 U118 ( .IN1(mem_data0[16]), .IN2(n2), .Q(N115) );
  AND2X1 U119 ( .IN1(mem_data0[15]), .IN2(n2), .Q(N114) );
  AND2X1 U120 ( .IN1(mem_data0[14]), .IN2(n2), .Q(N113) );
  AND2X1 U121 ( .IN1(mem_data0[13]), .IN2(n2), .Q(N112) );
  AND2X1 U122 ( .IN1(mem_data0[12]), .IN2(n2), .Q(N111) );
  AND2X1 U123 ( .IN1(mem_data0[11]), .IN2(n2), .Q(N110) );
  AND2X1 U124 ( .IN1(cur_pc0[8]), .IN2(n1), .Q(N11) );
  AND2X1 U125 ( .IN1(mem_data0[10]), .IN2(n1), .Q(N109) );
  AND2X1 U126 ( .IN1(mem_data0[9]), .IN2(n1), .Q(N108) );
  AND2X1 U127 ( .IN1(mem_data0[8]), .IN2(n1), .Q(N107) );
  AND2X1 U128 ( .IN1(mem_data0[7]), .IN2(n1), .Q(N106) );
  AND2X1 U129 ( .IN1(mem_data0[6]), .IN2(n1), .Q(N105) );
  AND2X1 U130 ( .IN1(mem_data0[5]), .IN2(n1), .Q(N104) );
  AND2X1 U131 ( .IN1(mem_data0[4]), .IN2(n1), .Q(N103) );
  AND2X1 U132 ( .IN1(mem_data0[3]), .IN2(n1), .Q(N102) );
  AND2X1 U133 ( .IN1(mem_data0[2]), .IN2(n1), .Q(N101) );
  AND2X1 U134 ( .IN1(mem_data0[1]), .IN2(n1), .Q(N100) );
  AND2X1 U135 ( .IN1(cur_pc0[7]), .IN2(n1), .Q(N10) );
  INVX0 U136 ( .INP(nrst), .ZN(n12) );
  INVX0 U137 ( .INP(n12), .ZN(n7) );
  INVX0 U138 ( .INP(n12), .ZN(n8) );
  INVX0 U139 ( .INP(n12), .ZN(n9) );
  INVX0 U140 ( .INP(n12), .ZN(n10) );
  INVX0 U141 ( .INP(n12), .ZN(n11) );
  INVX0 U142 ( .INP(n12), .ZN(n5) );
  INVX0 U143 ( .INP(n12), .ZN(n6) );
  INVX0 U144 ( .INP(n12), .ZN(n4) );
  INVX0 U145 ( .INP(n12), .ZN(n1) );
  INVX0 U146 ( .INP(n12), .ZN(n2) );
  INVX0 U147 ( .INP(n12), .ZN(n3) );
endmodule


module mem_wb_reg ( clk, nrst, cur_pc0, next_pc0, reg_data0, reg_addr0, cur_pc, 
        next_pc, reg_data, reg_addr );
  input [31:0] cur_pc0;
  input [31:0] next_pc0;
  input [31:0] reg_data0;
  input [4:0] reg_addr0;
  output [31:0] cur_pc;
  output [31:0] next_pc;
  output [31:0] reg_data;
  output [4:0] reg_addr;
  input clk, nrst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102;

  DFFX1 \reg_data_reg[31]  ( .D(N98), .CLK(clk), .Q(reg_data[31]) );
  DFFX1 \reg_data_reg[30]  ( .D(N97), .CLK(clk), .Q(reg_data[30]) );
  DFFX1 \reg_data_reg[29]  ( .D(N96), .CLK(clk), .Q(reg_data[29]) );
  DFFX1 \reg_data_reg[28]  ( .D(N95), .CLK(clk), .Q(reg_data[28]) );
  DFFX1 \reg_data_reg[27]  ( .D(N94), .CLK(clk), .Q(reg_data[27]) );
  DFFX1 \reg_data_reg[26]  ( .D(N93), .CLK(clk), .Q(reg_data[26]) );
  DFFX1 \reg_data_reg[25]  ( .D(N92), .CLK(clk), .Q(reg_data[25]) );
  DFFX1 \reg_data_reg[24]  ( .D(N91), .CLK(clk), .Q(reg_data[24]) );
  DFFX1 \reg_data_reg[23]  ( .D(N90), .CLK(clk), .Q(reg_data[23]) );
  DFFX1 \reg_data_reg[22]  ( .D(N89), .CLK(clk), .Q(reg_data[22]) );
  DFFX1 \reg_data_reg[21]  ( .D(N88), .CLK(clk), .Q(reg_data[21]) );
  DFFX1 \reg_data_reg[20]  ( .D(N87), .CLK(clk), .Q(reg_data[20]) );
  DFFX1 \reg_data_reg[19]  ( .D(N86), .CLK(clk), .Q(reg_data[19]) );
  DFFX1 \reg_data_reg[18]  ( .D(N85), .CLK(clk), .Q(reg_data[18]) );
  DFFX1 \reg_data_reg[17]  ( .D(N84), .CLK(clk), .Q(reg_data[17]) );
  DFFX1 \reg_data_reg[16]  ( .D(N83), .CLK(clk), .Q(reg_data[16]) );
  DFFX1 \reg_data_reg[15]  ( .D(N82), .CLK(clk), .Q(reg_data[15]) );
  DFFX1 \reg_data_reg[14]  ( .D(N81), .CLK(clk), .Q(reg_data[14]) );
  DFFX1 \reg_data_reg[13]  ( .D(N80), .CLK(clk), .Q(reg_data[13]) );
  DFFX1 \reg_data_reg[12]  ( .D(N79), .CLK(clk), .Q(reg_data[12]) );
  DFFX1 \reg_data_reg[11]  ( .D(N78), .CLK(clk), .Q(reg_data[11]) );
  DFFX1 \reg_data_reg[10]  ( .D(N77), .CLK(clk), .Q(reg_data[10]) );
  DFFX1 \reg_data_reg[9]  ( .D(N76), .CLK(clk), .Q(reg_data[9]) );
  DFFX1 \reg_data_reg[8]  ( .D(N75), .CLK(clk), .Q(reg_data[8]) );
  DFFX1 \reg_data_reg[7]  ( .D(N74), .CLK(clk), .Q(reg_data[7]) );
  DFFX1 \reg_data_reg[6]  ( .D(N73), .CLK(clk), .Q(reg_data[6]) );
  DFFX1 \reg_data_reg[5]  ( .D(N72), .CLK(clk), .Q(reg_data[5]) );
  DFFX1 \reg_data_reg[4]  ( .D(N71), .CLK(clk), .Q(reg_data[4]) );
  DFFX1 \reg_data_reg[3]  ( .D(N70), .CLK(clk), .Q(reg_data[3]) );
  DFFX1 \reg_data_reg[2]  ( .D(N69), .CLK(clk), .Q(reg_data[2]) );
  DFFX1 \reg_data_reg[1]  ( .D(N68), .CLK(clk), .Q(reg_data[1]) );
  DFFX1 \reg_data_reg[0]  ( .D(N67), .CLK(clk), .Q(reg_data[0]) );
  DFFX1 \reg_addr_reg[3]  ( .D(N102), .CLK(clk), .Q(reg_addr[3]) );
  DFFX1 \reg_addr_reg[2]  ( .D(N101), .CLK(clk), .Q(reg_addr[2]) );
  DFFX1 \reg_addr_reg[1]  ( .D(N100), .CLK(clk), .Q(reg_addr[1]) );
  DFFX1 \reg_addr_reg[0]  ( .D(N99), .CLK(clk), .Q(reg_addr[0]) );
  DFFX1 \cur_pc_reg[31]  ( .D(N34), .CLK(clk), .Q(cur_pc[31]) );
  DFFX1 \cur_pc_reg[30]  ( .D(N33), .CLK(clk), .Q(cur_pc[30]) );
  DFFX1 \cur_pc_reg[29]  ( .D(N32), .CLK(clk), .Q(cur_pc[29]) );
  DFFX1 \cur_pc_reg[28]  ( .D(N31), .CLK(clk), .Q(cur_pc[28]) );
  DFFX1 \cur_pc_reg[27]  ( .D(N30), .CLK(clk), .Q(cur_pc[27]) );
  DFFX1 \cur_pc_reg[26]  ( .D(N29), .CLK(clk), .Q(cur_pc[26]) );
  DFFX1 \cur_pc_reg[25]  ( .D(N28), .CLK(clk), .Q(cur_pc[25]) );
  DFFX1 \cur_pc_reg[24]  ( .D(N27), .CLK(clk), .Q(cur_pc[24]) );
  DFFX1 \cur_pc_reg[23]  ( .D(N26), .CLK(clk), .Q(cur_pc[23]) );
  DFFX1 \cur_pc_reg[22]  ( .D(N25), .CLK(clk), .Q(cur_pc[22]) );
  DFFX1 \cur_pc_reg[21]  ( .D(N24), .CLK(clk), .Q(cur_pc[21]) );
  DFFX1 \cur_pc_reg[20]  ( .D(N23), .CLK(clk), .Q(cur_pc[20]) );
  DFFX1 \cur_pc_reg[19]  ( .D(N22), .CLK(clk), .Q(cur_pc[19]) );
  DFFX1 \cur_pc_reg[18]  ( .D(N21), .CLK(clk), .Q(cur_pc[18]) );
  DFFX1 \cur_pc_reg[17]  ( .D(N20), .CLK(clk), .Q(cur_pc[17]) );
  DFFX1 \cur_pc_reg[16]  ( .D(N19), .CLK(clk), .Q(cur_pc[16]) );
  DFFX1 \cur_pc_reg[15]  ( .D(N18), .CLK(clk), .Q(cur_pc[15]) );
  DFFX1 \cur_pc_reg[14]  ( .D(N17), .CLK(clk), .Q(cur_pc[14]) );
  DFFX1 \cur_pc_reg[13]  ( .D(N16), .CLK(clk), .Q(cur_pc[13]) );
  DFFX1 \cur_pc_reg[12]  ( .D(N15), .CLK(clk), .Q(cur_pc[12]) );
  DFFX1 \cur_pc_reg[11]  ( .D(N14), .CLK(clk), .Q(cur_pc[11]) );
  DFFX1 \cur_pc_reg[10]  ( .D(N13), .CLK(clk), .Q(cur_pc[10]) );
  DFFX1 \cur_pc_reg[9]  ( .D(N12), .CLK(clk), .Q(cur_pc[9]) );
  DFFX1 \cur_pc_reg[8]  ( .D(N11), .CLK(clk), .Q(cur_pc[8]) );
  DFFX1 \cur_pc_reg[7]  ( .D(N10), .CLK(clk), .Q(cur_pc[7]) );
  DFFX1 \cur_pc_reg[6]  ( .D(N9), .CLK(clk), .Q(cur_pc[6]) );
  DFFX1 \cur_pc_reg[5]  ( .D(N8), .CLK(clk), .Q(cur_pc[5]) );
  DFFX1 \cur_pc_reg[4]  ( .D(N7), .CLK(clk), .Q(cur_pc[4]) );
  DFFX1 \cur_pc_reg[3]  ( .D(N6), .CLK(clk), .Q(cur_pc[3]) );
  DFFX1 \cur_pc_reg[2]  ( .D(N5), .CLK(clk), .Q(cur_pc[2]) );
  DFFX1 \cur_pc_reg[1]  ( .D(N4), .CLK(clk), .Q(cur_pc[1]) );
  DFFX1 \cur_pc_reg[0]  ( .D(N3), .CLK(clk), .Q(cur_pc[0]) );
  DFFX1 \next_pc_reg[31]  ( .D(N66), .CLK(clk), .Q(next_pc[31]) );
  DFFX1 \next_pc_reg[30]  ( .D(N65), .CLK(clk), .Q(next_pc[30]) );
  DFFX1 \next_pc_reg[29]  ( .D(N64), .CLK(clk), .Q(next_pc[29]) );
  DFFX1 \next_pc_reg[28]  ( .D(N63), .CLK(clk), .Q(next_pc[28]) );
  DFFX1 \next_pc_reg[27]  ( .D(N62), .CLK(clk), .Q(next_pc[27]) );
  DFFX1 \next_pc_reg[26]  ( .D(N61), .CLK(clk), .Q(next_pc[26]) );
  DFFX1 \next_pc_reg[25]  ( .D(N60), .CLK(clk), .Q(next_pc[25]) );
  DFFX1 \next_pc_reg[24]  ( .D(N59), .CLK(clk), .Q(next_pc[24]) );
  DFFX1 \next_pc_reg[23]  ( .D(N58), .CLK(clk), .Q(next_pc[23]) );
  DFFX1 \next_pc_reg[22]  ( .D(N57), .CLK(clk), .Q(next_pc[22]) );
  DFFX1 \next_pc_reg[21]  ( .D(N56), .CLK(clk), .Q(next_pc[21]) );
  DFFX1 \next_pc_reg[20]  ( .D(N55), .CLK(clk), .Q(next_pc[20]) );
  DFFX1 \next_pc_reg[19]  ( .D(N54), .CLK(clk), .Q(next_pc[19]) );
  DFFX1 \next_pc_reg[18]  ( .D(N53), .CLK(clk), .Q(next_pc[18]) );
  DFFX1 \next_pc_reg[17]  ( .D(N52), .CLK(clk), .Q(next_pc[17]) );
  DFFX1 \next_pc_reg[16]  ( .D(N51), .CLK(clk), .Q(next_pc[16]) );
  DFFX1 \next_pc_reg[15]  ( .D(N50), .CLK(clk), .Q(next_pc[15]) );
  DFFX1 \next_pc_reg[14]  ( .D(N49), .CLK(clk), .Q(next_pc[14]) );
  DFFX1 \next_pc_reg[13]  ( .D(N48), .CLK(clk), .Q(next_pc[13]) );
  DFFX1 \next_pc_reg[12]  ( .D(N47), .CLK(clk), .Q(next_pc[12]) );
  DFFX1 \next_pc_reg[11]  ( .D(N46), .CLK(clk), .Q(next_pc[11]) );
  DFFX1 \next_pc_reg[10]  ( .D(N45), .CLK(clk), .Q(next_pc[10]) );
  DFFX1 \next_pc_reg[9]  ( .D(N44), .CLK(clk), .Q(next_pc[9]) );
  DFFX1 \next_pc_reg[8]  ( .D(N43), .CLK(clk), .Q(next_pc[8]) );
  DFFX1 \next_pc_reg[7]  ( .D(N42), .CLK(clk), .Q(next_pc[7]) );
  DFFX1 \next_pc_reg[6]  ( .D(N41), .CLK(clk), .Q(next_pc[6]) );
  DFFX1 \next_pc_reg[5]  ( .D(N40), .CLK(clk), .Q(next_pc[5]) );
  DFFX1 \next_pc_reg[4]  ( .D(N39), .CLK(clk), .Q(next_pc[4]) );
  DFFX1 \next_pc_reg[3]  ( .D(N38), .CLK(clk), .Q(next_pc[3]) );
  DFFX1 \next_pc_reg[2]  ( .D(N37), .CLK(clk), .Q(next_pc[2]) );
  DFFX1 \next_pc_reg[1]  ( .D(N36), .CLK(clk), .Q(next_pc[1]) );
  DFFX1 \next_pc_reg[0]  ( .D(N35), .CLK(clk), .Q(next_pc[0]) );
  AND2X1 U3 ( .IN1(reg_addr0[0]), .IN2(nrst), .Q(N99) );
  AND2X1 U4 ( .IN1(reg_data0[31]), .IN2(nrst), .Q(N98) );
  AND2X1 U5 ( .IN1(reg_data0[30]), .IN2(nrst), .Q(N97) );
  AND2X1 U6 ( .IN1(reg_data0[29]), .IN2(nrst), .Q(N96) );
  AND2X1 U7 ( .IN1(reg_data0[28]), .IN2(nrst), .Q(N95) );
  AND2X1 U8 ( .IN1(reg_data0[27]), .IN2(nrst), .Q(N94) );
  AND2X1 U9 ( .IN1(reg_data0[26]), .IN2(nrst), .Q(N93) );
  AND2X1 U10 ( .IN1(reg_data0[25]), .IN2(nrst), .Q(N92) );
  AND2X1 U11 ( .IN1(reg_data0[24]), .IN2(nrst), .Q(N91) );
  AND2X1 U12 ( .IN1(reg_data0[23]), .IN2(nrst), .Q(N90) );
  AND2X1 U13 ( .IN1(cur_pc0[6]), .IN2(nrst), .Q(N9) );
  AND2X1 U14 ( .IN1(reg_data0[22]), .IN2(nrst), .Q(N89) );
  AND2X1 U15 ( .IN1(reg_data0[21]), .IN2(nrst), .Q(N88) );
  AND2X1 U16 ( .IN1(reg_data0[20]), .IN2(nrst), .Q(N87) );
  AND2X1 U17 ( .IN1(reg_data0[19]), .IN2(nrst), .Q(N86) );
  AND2X1 U18 ( .IN1(reg_data0[18]), .IN2(nrst), .Q(N85) );
  AND2X1 U19 ( .IN1(reg_data0[17]), .IN2(nrst), .Q(N84) );
  AND2X1 U20 ( .IN1(reg_data0[16]), .IN2(nrst), .Q(N83) );
  AND2X1 U21 ( .IN1(reg_data0[15]), .IN2(nrst), .Q(N82) );
  AND2X1 U22 ( .IN1(reg_data0[14]), .IN2(nrst), .Q(N81) );
  AND2X1 U23 ( .IN1(reg_data0[13]), .IN2(nrst), .Q(N80) );
  AND2X1 U24 ( .IN1(cur_pc0[5]), .IN2(nrst), .Q(N8) );
  AND2X1 U25 ( .IN1(reg_data0[12]), .IN2(nrst), .Q(N79) );
  AND2X1 U26 ( .IN1(reg_data0[11]), .IN2(nrst), .Q(N78) );
  AND2X1 U27 ( .IN1(reg_data0[10]), .IN2(nrst), .Q(N77) );
  AND2X1 U28 ( .IN1(reg_data0[9]), .IN2(nrst), .Q(N76) );
  AND2X1 U29 ( .IN1(reg_data0[8]), .IN2(nrst), .Q(N75) );
  AND2X1 U30 ( .IN1(reg_data0[7]), .IN2(nrst), .Q(N74) );
  AND2X1 U31 ( .IN1(reg_data0[6]), .IN2(nrst), .Q(N73) );
  AND2X1 U32 ( .IN1(reg_data0[5]), .IN2(nrst), .Q(N72) );
  AND2X1 U33 ( .IN1(reg_data0[4]), .IN2(nrst), .Q(N71) );
  AND2X1 U34 ( .IN1(reg_data0[3]), .IN2(nrst), .Q(N70) );
  AND2X1 U35 ( .IN1(cur_pc0[4]), .IN2(nrst), .Q(N7) );
  AND2X1 U36 ( .IN1(reg_data0[2]), .IN2(nrst), .Q(N69) );
  AND2X1 U37 ( .IN1(reg_data0[1]), .IN2(nrst), .Q(N68) );
  AND2X1 U38 ( .IN1(reg_data0[0]), .IN2(nrst), .Q(N67) );
  AND2X1 U39 ( .IN1(next_pc0[31]), .IN2(nrst), .Q(N66) );
  AND2X1 U40 ( .IN1(next_pc0[30]), .IN2(nrst), .Q(N65) );
  AND2X1 U41 ( .IN1(next_pc0[29]), .IN2(nrst), .Q(N64) );
  AND2X1 U42 ( .IN1(next_pc0[28]), .IN2(nrst), .Q(N63) );
  AND2X1 U43 ( .IN1(next_pc0[27]), .IN2(nrst), .Q(N62) );
  AND2X1 U44 ( .IN1(next_pc0[26]), .IN2(nrst), .Q(N61) );
  AND2X1 U45 ( .IN1(next_pc0[25]), .IN2(nrst), .Q(N60) );
  AND2X1 U46 ( .IN1(cur_pc0[3]), .IN2(nrst), .Q(N6) );
  AND2X1 U47 ( .IN1(next_pc0[24]), .IN2(nrst), .Q(N59) );
  AND2X1 U48 ( .IN1(next_pc0[23]), .IN2(nrst), .Q(N58) );
  AND2X1 U49 ( .IN1(next_pc0[22]), .IN2(nrst), .Q(N57) );
  AND2X1 U50 ( .IN1(next_pc0[21]), .IN2(nrst), .Q(N56) );
  AND2X1 U51 ( .IN1(next_pc0[20]), .IN2(nrst), .Q(N55) );
  AND2X1 U52 ( .IN1(next_pc0[19]), .IN2(nrst), .Q(N54) );
  AND2X1 U53 ( .IN1(next_pc0[18]), .IN2(nrst), .Q(N53) );
  AND2X1 U54 ( .IN1(next_pc0[17]), .IN2(nrst), .Q(N52) );
  AND2X1 U55 ( .IN1(next_pc0[16]), .IN2(nrst), .Q(N51) );
  AND2X1 U56 ( .IN1(next_pc0[15]), .IN2(nrst), .Q(N50) );
  AND2X1 U57 ( .IN1(cur_pc0[2]), .IN2(nrst), .Q(N5) );
  AND2X1 U58 ( .IN1(next_pc0[14]), .IN2(nrst), .Q(N49) );
  AND2X1 U59 ( .IN1(next_pc0[13]), .IN2(nrst), .Q(N48) );
  AND2X1 U60 ( .IN1(next_pc0[12]), .IN2(nrst), .Q(N47) );
  AND2X1 U61 ( .IN1(next_pc0[11]), .IN2(nrst), .Q(N46) );
  AND2X1 U62 ( .IN1(next_pc0[10]), .IN2(nrst), .Q(N45) );
  AND2X1 U63 ( .IN1(next_pc0[9]), .IN2(nrst), .Q(N44) );
  AND2X1 U64 ( .IN1(next_pc0[8]), .IN2(nrst), .Q(N43) );
  AND2X1 U65 ( .IN1(next_pc0[7]), .IN2(nrst), .Q(N42) );
  AND2X1 U66 ( .IN1(next_pc0[6]), .IN2(nrst), .Q(N41) );
  AND2X1 U67 ( .IN1(next_pc0[5]), .IN2(nrst), .Q(N40) );
  AND2X1 U68 ( .IN1(cur_pc0[1]), .IN2(nrst), .Q(N4) );
  AND2X1 U69 ( .IN1(next_pc0[4]), .IN2(nrst), .Q(N39) );
  AND2X1 U70 ( .IN1(next_pc0[3]), .IN2(nrst), .Q(N38) );
  AND2X1 U71 ( .IN1(next_pc0[2]), .IN2(nrst), .Q(N37) );
  AND2X1 U72 ( .IN1(next_pc0[1]), .IN2(nrst), .Q(N36) );
  AND2X1 U73 ( .IN1(next_pc0[0]), .IN2(nrst), .Q(N35) );
  AND2X1 U74 ( .IN1(cur_pc0[31]), .IN2(nrst), .Q(N34) );
  AND2X1 U75 ( .IN1(cur_pc0[30]), .IN2(nrst), .Q(N33) );
  AND2X1 U76 ( .IN1(cur_pc0[29]), .IN2(nrst), .Q(N32) );
  AND2X1 U77 ( .IN1(cur_pc0[28]), .IN2(nrst), .Q(N31) );
  AND2X1 U78 ( .IN1(cur_pc0[27]), .IN2(nrst), .Q(N30) );
  AND2X1 U79 ( .IN1(cur_pc0[0]), .IN2(nrst), .Q(N3) );
  AND2X1 U80 ( .IN1(cur_pc0[26]), .IN2(nrst), .Q(N29) );
  AND2X1 U81 ( .IN1(cur_pc0[25]), .IN2(nrst), .Q(N28) );
  AND2X1 U82 ( .IN1(cur_pc0[24]), .IN2(nrst), .Q(N27) );
  AND2X1 U83 ( .IN1(cur_pc0[23]), .IN2(nrst), .Q(N26) );
  AND2X1 U84 ( .IN1(cur_pc0[22]), .IN2(nrst), .Q(N25) );
  AND2X1 U85 ( .IN1(cur_pc0[21]), .IN2(nrst), .Q(N24) );
  AND2X1 U86 ( .IN1(cur_pc0[20]), .IN2(nrst), .Q(N23) );
  AND2X1 U87 ( .IN1(cur_pc0[19]), .IN2(nrst), .Q(N22) );
  AND2X1 U88 ( .IN1(cur_pc0[18]), .IN2(nrst), .Q(N21) );
  AND2X1 U89 ( .IN1(cur_pc0[17]), .IN2(nrst), .Q(N20) );
  AND2X1 U90 ( .IN1(cur_pc0[16]), .IN2(nrst), .Q(N19) );
  AND2X1 U91 ( .IN1(cur_pc0[15]), .IN2(nrst), .Q(N18) );
  AND2X1 U92 ( .IN1(cur_pc0[14]), .IN2(nrst), .Q(N17) );
  AND2X1 U93 ( .IN1(cur_pc0[13]), .IN2(nrst), .Q(N16) );
  AND2X1 U94 ( .IN1(cur_pc0[12]), .IN2(nrst), .Q(N15) );
  AND2X1 U95 ( .IN1(cur_pc0[11]), .IN2(nrst), .Q(N14) );
  AND2X1 U96 ( .IN1(cur_pc0[10]), .IN2(nrst), .Q(N13) );
  AND2X1 U97 ( .IN1(cur_pc0[9]), .IN2(nrst), .Q(N12) );
  AND2X1 U98 ( .IN1(cur_pc0[8]), .IN2(nrst), .Q(N11) );
  AND2X1 U100 ( .IN1(reg_addr0[3]), .IN2(nrst), .Q(N102) );
  AND2X1 U101 ( .IN1(reg_addr0[2]), .IN2(nrst), .Q(N101) );
  AND2X1 U102 ( .IN1(reg_addr0[1]), .IN2(nrst), .Q(N100) );
  AND2X1 U103 ( .IN1(cur_pc0[7]), .IN2(nrst), .Q(N10) );
  DFFSSRX1 \reg_addr_reg[4]  ( .D(reg_addr0[4]), .RSTB(nrst), .SETB(1'b1), 
        .CLK(clk), .Q(reg_addr[4]) );
endmodule


module reg32_5 ( clk, nrst, en, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, nrst, en;
  wire   n1, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69;

  DFFX1 \data_out_reg[31]  ( .D(n36), .CLK(clk), .Q(data_out[31]) );
  DFFX1 \data_out_reg[30]  ( .D(n37), .CLK(clk), .Q(data_out[30]) );
  DFFX1 \data_out_reg[29]  ( .D(n38), .CLK(clk), .Q(data_out[29]) );
  DFFX1 \data_out_reg[28]  ( .D(n39), .CLK(clk), .Q(data_out[28]) );
  DFFX1 \data_out_reg[27]  ( .D(n40), .CLK(clk), .Q(data_out[27]) );
  DFFX1 \data_out_reg[26]  ( .D(n41), .CLK(clk), .Q(data_out[26]) );
  DFFX1 \data_out_reg[25]  ( .D(n42), .CLK(clk), .Q(data_out[25]) );
  DFFX1 \data_out_reg[24]  ( .D(n43), .CLK(clk), .Q(data_out[24]) );
  DFFX1 \data_out_reg[23]  ( .D(n44), .CLK(clk), .Q(data_out[23]) );
  DFFX1 \data_out_reg[22]  ( .D(n45), .CLK(clk), .Q(data_out[22]) );
  DFFX1 \data_out_reg[21]  ( .D(n46), .CLK(clk), .Q(data_out[21]) );
  DFFX1 \data_out_reg[20]  ( .D(n47), .CLK(clk), .Q(data_out[20]) );
  DFFX1 \data_out_reg[19]  ( .D(n48), .CLK(clk), .Q(data_out[19]) );
  DFFX1 \data_out_reg[18]  ( .D(n49), .CLK(clk), .Q(data_out[18]) );
  DFFX1 \data_out_reg[17]  ( .D(n50), .CLK(clk), .Q(data_out[17]) );
  DFFX1 \data_out_reg[16]  ( .D(n51), .CLK(clk), .Q(data_out[16]) );
  DFFX1 \data_out_reg[15]  ( .D(n52), .CLK(clk), .Q(data_out[15]) );
  DFFX1 \data_out_reg[14]  ( .D(n53), .CLK(clk), .Q(data_out[14]) );
  DFFX1 \data_out_reg[13]  ( .D(n54), .CLK(clk), .Q(data_out[13]) );
  DFFX1 \data_out_reg[12]  ( .D(n55), .CLK(clk), .Q(data_out[12]) );
  DFFX1 \data_out_reg[11]  ( .D(n56), .CLK(clk), .Q(data_out[11]) );
  DFFX1 \data_out_reg[10]  ( .D(n57), .CLK(clk), .Q(data_out[10]) );
  DFFX1 \data_out_reg[9]  ( .D(n58), .CLK(clk), .Q(data_out[9]) );
  DFFX1 \data_out_reg[8]  ( .D(n59), .CLK(clk), .Q(data_out[8]) );
  DFFX1 \data_out_reg[7]  ( .D(n60), .CLK(clk), .Q(data_out[7]) );
  DFFX1 \data_out_reg[6]  ( .D(n61), .CLK(clk), .Q(data_out[6]) );
  DFFX1 \data_out_reg[5]  ( .D(n62), .CLK(clk), .Q(data_out[5]) );
  DFFX1 \data_out_reg[4]  ( .D(n63), .CLK(clk), .Q(data_out[4]) );
  DFFX1 \data_out_reg[3]  ( .D(n64), .CLK(clk), .Q(data_out[3]) );
  DFFX1 \data_out_reg[2]  ( .D(n65), .CLK(clk), .Q(data_out[2]) );
  DFFX1 \data_out_reg[1]  ( .D(n66), .CLK(clk), .Q(data_out[1]) );
  DFFX1 \data_out_reg[0]  ( .D(n67), .CLK(clk), .Q(data_out[0]) );
  AO22X1 U4 ( .IN1(data_out[0]), .IN2(n69), .IN3(data_in[0]), .IN4(n1), .Q(n67) );
  AO22X1 U5 ( .IN1(data_out[1]), .IN2(n69), .IN3(data_in[1]), .IN4(n1), .Q(n66) );
  AO22X1 U6 ( .IN1(data_out[2]), .IN2(n69), .IN3(data_in[2]), .IN4(n1), .Q(n65) );
  AO22X1 U7 ( .IN1(data_out[3]), .IN2(n69), .IN3(data_in[3]), .IN4(n1), .Q(n64) );
  AO22X1 U8 ( .IN1(data_out[4]), .IN2(n69), .IN3(data_in[4]), .IN4(n1), .Q(n63) );
  AO22X1 U9 ( .IN1(data_out[5]), .IN2(n69), .IN3(data_in[5]), .IN4(n1), .Q(n62) );
  AO22X1 U10 ( .IN1(data_out[6]), .IN2(n69), .IN3(data_in[6]), .IN4(n1), .Q(
        n61) );
  AO22X1 U11 ( .IN1(data_out[7]), .IN2(n69), .IN3(data_in[7]), .IN4(n1), .Q(
        n60) );
  AO22X1 U12 ( .IN1(data_out[8]), .IN2(n69), .IN3(data_in[8]), .IN4(n1), .Q(
        n59) );
  AO22X1 U13 ( .IN1(data_out[9]), .IN2(n69), .IN3(data_in[9]), .IN4(n1), .Q(
        n58) );
  AO22X1 U14 ( .IN1(data_out[10]), .IN2(n69), .IN3(data_in[10]), .IN4(n1), .Q(
        n57) );
  AO22X1 U15 ( .IN1(data_out[11]), .IN2(n69), .IN3(data_in[11]), .IN4(n1), .Q(
        n56) );
  AO22X1 U16 ( .IN1(data_out[12]), .IN2(n69), .IN3(data_in[12]), .IN4(n1), .Q(
        n55) );
  AO22X1 U17 ( .IN1(data_out[13]), .IN2(n69), .IN3(data_in[13]), .IN4(n1), .Q(
        n54) );
  AO22X1 U18 ( .IN1(data_out[14]), .IN2(n69), .IN3(data_in[14]), .IN4(n1), .Q(
        n53) );
  AO22X1 U19 ( .IN1(data_out[15]), .IN2(n69), .IN3(data_in[15]), .IN4(n1), .Q(
        n52) );
  AO22X1 U20 ( .IN1(data_out[16]), .IN2(n69), .IN3(data_in[16]), .IN4(n1), .Q(
        n51) );
  AO22X1 U21 ( .IN1(data_out[17]), .IN2(n69), .IN3(data_in[17]), .IN4(n1), .Q(
        n50) );
  AO22X1 U22 ( .IN1(data_out[18]), .IN2(n69), .IN3(data_in[18]), .IN4(n1), .Q(
        n49) );
  AO22X1 U23 ( .IN1(data_out[19]), .IN2(n69), .IN3(data_in[19]), .IN4(n1), .Q(
        n48) );
  AO22X1 U24 ( .IN1(data_out[20]), .IN2(n69), .IN3(data_in[20]), .IN4(n1), .Q(
        n47) );
  AO22X1 U25 ( .IN1(data_out[21]), .IN2(n69), .IN3(data_in[21]), .IN4(n1), .Q(
        n46) );
  AO22X1 U26 ( .IN1(data_out[22]), .IN2(n69), .IN3(data_in[22]), .IN4(n1), .Q(
        n45) );
  AO22X1 U27 ( .IN1(data_out[23]), .IN2(n69), .IN3(data_in[23]), .IN4(n1), .Q(
        n44) );
  AO22X1 U28 ( .IN1(data_out[24]), .IN2(n69), .IN3(data_in[24]), .IN4(n1), .Q(
        n43) );
  AO22X1 U29 ( .IN1(data_out[25]), .IN2(n69), .IN3(data_in[25]), .IN4(n1), .Q(
        n42) );
  AO22X1 U30 ( .IN1(data_out[26]), .IN2(n69), .IN3(data_in[26]), .IN4(n1), .Q(
        n41) );
  AO22X1 U31 ( .IN1(data_out[27]), .IN2(n69), .IN3(data_in[27]), .IN4(n1), .Q(
        n40) );
  AO22X1 U32 ( .IN1(data_out[28]), .IN2(n69), .IN3(data_in[28]), .IN4(n1), .Q(
        n39) );
  AO22X1 U33 ( .IN1(data_out[29]), .IN2(n69), .IN3(data_in[29]), .IN4(n1), .Q(
        n38) );
  AO22X1 U34 ( .IN1(data_out[30]), .IN2(n69), .IN3(data_in[30]), .IN4(n1), .Q(
        n37) );
  AO22X1 U35 ( .IN1(data_out[31]), .IN2(n69), .IN3(data_in[31]), .IN4(n1), .Q(
        n36) );
  INVX0 U2 ( .INP(n68), .ZN(n1) );
  AND2X1 U3 ( .IN1(nrst), .IN2(n68), .Q(n69) );
  NAND2X1 U36 ( .IN1(nrst), .IN2(en), .QN(n68) );
endmodule


module reg_fwd ( clk, nrst, fwd_opA0, fwd_opB0, fwd_jr0, fwd_opA, fwd_opB, 
        fwd_sw, fwd_jr );
  input [2:0] fwd_opA0;
  input [2:0] fwd_opB0;
  input [2:0] fwd_jr0;
  output [2:0] fwd_opA;
  output [2:0] fwd_opB;
  output [2:0] fwd_sw;
  output [2:0] fwd_jr;
  input clk, nrst;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11;
  assign fwd_jr[2] = fwd_jr0[2];
  assign fwd_jr[1] = fwd_jr0[1];
  assign fwd_jr[0] = fwd_jr0[0];

  DFFX1 \fwd_opB_reg[2]  ( .D(N8), .CLK(clk), .Q(fwd_opB[2]) );
  DFFX1 \fwd_opB_reg[1]  ( .D(N7), .CLK(clk), .Q(fwd_opB[1]) );
  DFFX1 \fwd_opB_reg[0]  ( .D(N6), .CLK(clk), .Q(fwd_opB[0]) );
  DFFX1 \fwd_sw_reg[2]  ( .D(N11), .CLK(clk), .Q(fwd_sw[2]) );
  DFFX1 \fwd_sw_reg[1]  ( .D(N10), .CLK(clk), .Q(fwd_sw[1]) );
  DFFX1 \fwd_sw_reg[0]  ( .D(N9), .CLK(clk), .Q(fwd_sw[0]) );
  DFFX1 \fwd_opA_reg[2]  ( .D(N5), .CLK(clk), .Q(fwd_opA[2]) );
  DFFX1 \fwd_opA_reg[1]  ( .D(N4), .CLK(clk), .Q(fwd_opA[1]) );
  DFFX1 \fwd_opA_reg[0]  ( .D(N3), .CLK(clk), .Q(fwd_opA[0]) );
  AND2X1 U3 ( .IN1(nrst), .IN2(fwd_jr0[0]), .Q(N9) );
  AND2X1 U4 ( .IN1(fwd_opB0[2]), .IN2(nrst), .Q(N8) );
  AND2X1 U5 ( .IN1(fwd_opB0[1]), .IN2(nrst), .Q(N7) );
  AND2X1 U6 ( .IN1(fwd_opB0[0]), .IN2(nrst), .Q(N6) );
  AND2X1 U7 ( .IN1(fwd_opA0[2]), .IN2(nrst), .Q(N5) );
  AND2X1 U8 ( .IN1(fwd_opA0[1]), .IN2(nrst), .Q(N4) );
  AND2X1 U9 ( .IN1(fwd_opA0[0]), .IN2(nrst), .Q(N3) );
  AND2X1 U10 ( .IN1(fwd_jr0[2]), .IN2(nrst), .Q(N11) );
  AND2X1 U11 ( .IN1(fwd_jr0[1]), .IN2(nrst), .Q(N10) );
endmodule


module reg32_4 ( clk, nrst, en, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, nrst, en;
  wire   n1, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70;

  DFFX1 \data_out_reg[31]  ( .D(n37), .CLK(clk), .Q(data_out[31]) );
  DFFX1 \data_out_reg[30]  ( .D(n38), .CLK(clk), .Q(data_out[30]) );
  DFFX1 \data_out_reg[29]  ( .D(n39), .CLK(clk), .Q(data_out[29]) );
  DFFX1 \data_out_reg[28]  ( .D(n40), .CLK(clk), .Q(data_out[28]) );
  DFFX1 \data_out_reg[27]  ( .D(n41), .CLK(clk), .Q(data_out[27]) );
  DFFX1 \data_out_reg[26]  ( .D(n42), .CLK(clk), .Q(data_out[26]) );
  DFFX1 \data_out_reg[25]  ( .D(n43), .CLK(clk), .Q(data_out[25]) );
  DFFX1 \data_out_reg[24]  ( .D(n44), .CLK(clk), .Q(data_out[24]) );
  DFFX1 \data_out_reg[23]  ( .D(n45), .CLK(clk), .Q(data_out[23]) );
  DFFX1 \data_out_reg[22]  ( .D(n46), .CLK(clk), .Q(data_out[22]) );
  DFFX1 \data_out_reg[21]  ( .D(n47), .CLK(clk), .Q(data_out[21]) );
  DFFX1 \data_out_reg[20]  ( .D(n48), .CLK(clk), .Q(data_out[20]) );
  DFFX1 \data_out_reg[19]  ( .D(n49), .CLK(clk), .Q(data_out[19]) );
  DFFX1 \data_out_reg[18]  ( .D(n50), .CLK(clk), .Q(data_out[18]) );
  DFFX1 \data_out_reg[17]  ( .D(n51), .CLK(clk), .Q(data_out[17]) );
  DFFX1 \data_out_reg[16]  ( .D(n52), .CLK(clk), .Q(data_out[16]) );
  DFFX1 \data_out_reg[15]  ( .D(n53), .CLK(clk), .Q(data_out[15]) );
  DFFX1 \data_out_reg[14]  ( .D(n54), .CLK(clk), .Q(data_out[14]) );
  DFFX1 \data_out_reg[13]  ( .D(n55), .CLK(clk), .Q(data_out[13]) );
  DFFX1 \data_out_reg[12]  ( .D(n56), .CLK(clk), .Q(data_out[12]) );
  DFFX1 \data_out_reg[11]  ( .D(n57), .CLK(clk), .Q(data_out[11]) );
  DFFX1 \data_out_reg[10]  ( .D(n58), .CLK(clk), .Q(data_out[10]) );
  DFFX1 \data_out_reg[9]  ( .D(n59), .CLK(clk), .Q(data_out[9]) );
  DFFX1 \data_out_reg[8]  ( .D(n60), .CLK(clk), .Q(data_out[8]) );
  DFFX1 \data_out_reg[7]  ( .D(n61), .CLK(clk), .Q(data_out[7]) );
  DFFX1 \data_out_reg[6]  ( .D(n62), .CLK(clk), .Q(data_out[6]) );
  DFFX1 \data_out_reg[5]  ( .D(n63), .CLK(clk), .Q(data_out[5]) );
  DFFX1 \data_out_reg[4]  ( .D(n64), .CLK(clk), .Q(data_out[4]) );
  DFFX1 \data_out_reg[3]  ( .D(n65), .CLK(clk), .Q(data_out[3]) );
  DFFX1 \data_out_reg[2]  ( .D(n66), .CLK(clk), .Q(data_out[2]) );
  DFFX1 \data_out_reg[1]  ( .D(n67), .CLK(clk), .Q(data_out[1]) );
  DFFX1 \data_out_reg[0]  ( .D(n68), .CLK(clk), .Q(data_out[0]) );
  AO22X1 U4 ( .IN1(data_out[0]), .IN2(n70), .IN3(data_in[0]), .IN4(n36), .Q(
        n68) );
  AO22X1 U5 ( .IN1(data_out[1]), .IN2(n1), .IN3(data_in[1]), .IN4(n36), .Q(n67) );
  AO22X1 U6 ( .IN1(data_out[2]), .IN2(n70), .IN3(data_in[2]), .IN4(n36), .Q(
        n66) );
  AO22X1 U7 ( .IN1(data_out[3]), .IN2(n1), .IN3(data_in[3]), .IN4(n36), .Q(n65) );
  AO22X1 U8 ( .IN1(data_out[4]), .IN2(n70), .IN3(data_in[4]), .IN4(n36), .Q(
        n64) );
  AO22X1 U9 ( .IN1(data_out[5]), .IN2(n1), .IN3(data_in[5]), .IN4(n36), .Q(n63) );
  AO22X1 U10 ( .IN1(data_out[6]), .IN2(n70), .IN3(data_in[6]), .IN4(n36), .Q(
        n62) );
  AO22X1 U11 ( .IN1(data_out[7]), .IN2(n1), .IN3(data_in[7]), .IN4(n36), .Q(
        n61) );
  AO22X1 U12 ( .IN1(data_out[8]), .IN2(n70), .IN3(data_in[8]), .IN4(n36), .Q(
        n60) );
  AO22X1 U13 ( .IN1(data_out[9]), .IN2(n1), .IN3(data_in[9]), .IN4(n36), .Q(
        n59) );
  AO22X1 U14 ( .IN1(data_out[10]), .IN2(n70), .IN3(data_in[10]), .IN4(n36), 
        .Q(n58) );
  AO22X1 U15 ( .IN1(data_out[11]), .IN2(n1), .IN3(data_in[11]), .IN4(n36), .Q(
        n57) );
  AO22X1 U16 ( .IN1(data_out[12]), .IN2(n70), .IN3(data_in[12]), .IN4(n36), 
        .Q(n56) );
  AO22X1 U17 ( .IN1(data_out[13]), .IN2(n1), .IN3(data_in[13]), .IN4(n36), .Q(
        n55) );
  AO22X1 U18 ( .IN1(data_out[14]), .IN2(n70), .IN3(data_in[14]), .IN4(n36), 
        .Q(n54) );
  AO22X1 U19 ( .IN1(data_out[15]), .IN2(n1), .IN3(data_in[15]), .IN4(n36), .Q(
        n53) );
  AO22X1 U20 ( .IN1(data_out[16]), .IN2(n70), .IN3(data_in[16]), .IN4(n36), 
        .Q(n52) );
  AO22X1 U21 ( .IN1(data_out[17]), .IN2(n1), .IN3(data_in[17]), .IN4(n36), .Q(
        n51) );
  AO22X1 U22 ( .IN1(data_out[18]), .IN2(n70), .IN3(data_in[18]), .IN4(n36), 
        .Q(n50) );
  AO22X1 U23 ( .IN1(data_out[19]), .IN2(n1), .IN3(data_in[19]), .IN4(n36), .Q(
        n49) );
  AO22X1 U24 ( .IN1(data_out[20]), .IN2(n70), .IN3(data_in[20]), .IN4(n36), 
        .Q(n48) );
  AO22X1 U25 ( .IN1(data_out[21]), .IN2(n1), .IN3(data_in[21]), .IN4(n36), .Q(
        n47) );
  AO22X1 U26 ( .IN1(data_out[22]), .IN2(n70), .IN3(data_in[22]), .IN4(n36), 
        .Q(n46) );
  AO22X1 U27 ( .IN1(data_out[23]), .IN2(n1), .IN3(data_in[23]), .IN4(n36), .Q(
        n45) );
  AO22X1 U28 ( .IN1(data_out[24]), .IN2(n70), .IN3(data_in[24]), .IN4(n36), 
        .Q(n44) );
  AO22X1 U29 ( .IN1(data_out[25]), .IN2(n1), .IN3(data_in[25]), .IN4(n36), .Q(
        n43) );
  AO22X1 U30 ( .IN1(data_out[26]), .IN2(n70), .IN3(data_in[26]), .IN4(n36), 
        .Q(n42) );
  AO22X1 U31 ( .IN1(data_out[27]), .IN2(n1), .IN3(data_in[27]), .IN4(n36), .Q(
        n41) );
  AO22X1 U32 ( .IN1(data_out[28]), .IN2(n70), .IN3(data_in[28]), .IN4(n36), 
        .Q(n40) );
  AO22X1 U33 ( .IN1(data_out[29]), .IN2(n1), .IN3(data_in[29]), .IN4(n36), .Q(
        n39) );
  AO22X1 U34 ( .IN1(data_out[30]), .IN2(n70), .IN3(data_in[30]), .IN4(n36), 
        .Q(n38) );
  AO22X1 U35 ( .IN1(data_out[31]), .IN2(n1), .IN3(data_in[31]), .IN4(n36), .Q(
        n37) );
  INVX0 U2 ( .INP(n69), .ZN(n36) );
  AND2X1 U3 ( .IN1(nrst), .IN2(n69), .Q(n70) );
  AND2X1 U36 ( .IN1(nrst), .IN2(n69), .Q(n1) );
  NAND2X1 U37 ( .IN1(nrst), .IN2(en), .QN(n69) );
endmodule


module reg32_3 ( clk, nrst, en, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, nrst, en;
  wire   n1, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70;

  DFFX1 \data_out_reg[31]  ( .D(n37), .CLK(clk), .Q(data_out[31]) );
  DFFX1 \data_out_reg[30]  ( .D(n38), .CLK(clk), .Q(data_out[30]) );
  DFFX1 \data_out_reg[29]  ( .D(n39), .CLK(clk), .Q(data_out[29]) );
  DFFX1 \data_out_reg[28]  ( .D(n40), .CLK(clk), .Q(data_out[28]) );
  DFFX1 \data_out_reg[27]  ( .D(n41), .CLK(clk), .Q(data_out[27]) );
  DFFX1 \data_out_reg[26]  ( .D(n42), .CLK(clk), .Q(data_out[26]) );
  DFFX1 \data_out_reg[25]  ( .D(n43), .CLK(clk), .Q(data_out[25]) );
  DFFX1 \data_out_reg[24]  ( .D(n44), .CLK(clk), .Q(data_out[24]) );
  DFFX1 \data_out_reg[23]  ( .D(n45), .CLK(clk), .Q(data_out[23]) );
  DFFX1 \data_out_reg[22]  ( .D(n46), .CLK(clk), .Q(data_out[22]) );
  DFFX1 \data_out_reg[21]  ( .D(n47), .CLK(clk), .Q(data_out[21]) );
  DFFX1 \data_out_reg[20]  ( .D(n48), .CLK(clk), .Q(data_out[20]) );
  DFFX1 \data_out_reg[19]  ( .D(n49), .CLK(clk), .Q(data_out[19]) );
  DFFX1 \data_out_reg[18]  ( .D(n50), .CLK(clk), .Q(data_out[18]) );
  DFFX1 \data_out_reg[17]  ( .D(n51), .CLK(clk), .Q(data_out[17]) );
  DFFX1 \data_out_reg[16]  ( .D(n52), .CLK(clk), .Q(data_out[16]) );
  DFFX1 \data_out_reg[15]  ( .D(n53), .CLK(clk), .Q(data_out[15]) );
  DFFX1 \data_out_reg[14]  ( .D(n54), .CLK(clk), .Q(data_out[14]) );
  DFFX1 \data_out_reg[13]  ( .D(n55), .CLK(clk), .Q(data_out[13]) );
  DFFX1 \data_out_reg[12]  ( .D(n56), .CLK(clk), .Q(data_out[12]) );
  DFFX1 \data_out_reg[11]  ( .D(n57), .CLK(clk), .Q(data_out[11]) );
  DFFX1 \data_out_reg[10]  ( .D(n58), .CLK(clk), .Q(data_out[10]) );
  DFFX1 \data_out_reg[9]  ( .D(n59), .CLK(clk), .Q(data_out[9]) );
  DFFX1 \data_out_reg[8]  ( .D(n60), .CLK(clk), .Q(data_out[8]) );
  DFFX1 \data_out_reg[7]  ( .D(n61), .CLK(clk), .Q(data_out[7]) );
  DFFX1 \data_out_reg[6]  ( .D(n62), .CLK(clk), .Q(data_out[6]) );
  DFFX1 \data_out_reg[5]  ( .D(n63), .CLK(clk), .Q(data_out[5]) );
  DFFX1 \data_out_reg[4]  ( .D(n64), .CLK(clk), .Q(data_out[4]) );
  DFFX1 \data_out_reg[3]  ( .D(n65), .CLK(clk), .Q(data_out[3]) );
  DFFX1 \data_out_reg[2]  ( .D(n66), .CLK(clk), .Q(data_out[2]) );
  DFFX1 \data_out_reg[1]  ( .D(n67), .CLK(clk), .Q(data_out[1]) );
  DFFX1 \data_out_reg[0]  ( .D(n68), .CLK(clk), .Q(data_out[0]) );
  AO22X1 U4 ( .IN1(data_out[0]), .IN2(n70), .IN3(data_in[0]), .IN4(n36), .Q(
        n68) );
  AO22X1 U5 ( .IN1(data_out[1]), .IN2(n1), .IN3(data_in[1]), .IN4(n36), .Q(n67) );
  AO22X1 U6 ( .IN1(data_out[2]), .IN2(n70), .IN3(data_in[2]), .IN4(n36), .Q(
        n66) );
  AO22X1 U7 ( .IN1(data_out[3]), .IN2(n1), .IN3(data_in[3]), .IN4(n36), .Q(n65) );
  AO22X1 U8 ( .IN1(data_out[4]), .IN2(n70), .IN3(data_in[4]), .IN4(n36), .Q(
        n64) );
  AO22X1 U9 ( .IN1(data_out[5]), .IN2(n1), .IN3(data_in[5]), .IN4(n36), .Q(n63) );
  AO22X1 U10 ( .IN1(data_out[6]), .IN2(n70), .IN3(data_in[6]), .IN4(n36), .Q(
        n62) );
  AO22X1 U11 ( .IN1(data_out[7]), .IN2(n1), .IN3(data_in[7]), .IN4(n36), .Q(
        n61) );
  AO22X1 U12 ( .IN1(data_out[8]), .IN2(n70), .IN3(data_in[8]), .IN4(n36), .Q(
        n60) );
  AO22X1 U13 ( .IN1(data_out[9]), .IN2(n1), .IN3(data_in[9]), .IN4(n36), .Q(
        n59) );
  AO22X1 U14 ( .IN1(data_out[10]), .IN2(n70), .IN3(data_in[10]), .IN4(n36), 
        .Q(n58) );
  AO22X1 U15 ( .IN1(data_out[11]), .IN2(n1), .IN3(data_in[11]), .IN4(n36), .Q(
        n57) );
  AO22X1 U16 ( .IN1(data_out[12]), .IN2(n70), .IN3(data_in[12]), .IN4(n36), 
        .Q(n56) );
  AO22X1 U17 ( .IN1(data_out[13]), .IN2(n1), .IN3(data_in[13]), .IN4(n36), .Q(
        n55) );
  AO22X1 U18 ( .IN1(data_out[14]), .IN2(n70), .IN3(data_in[14]), .IN4(n36), 
        .Q(n54) );
  AO22X1 U19 ( .IN1(data_out[15]), .IN2(n1), .IN3(data_in[15]), .IN4(n36), .Q(
        n53) );
  AO22X1 U20 ( .IN1(data_out[16]), .IN2(n70), .IN3(data_in[16]), .IN4(n36), 
        .Q(n52) );
  AO22X1 U21 ( .IN1(data_out[17]), .IN2(n1), .IN3(data_in[17]), .IN4(n36), .Q(
        n51) );
  AO22X1 U22 ( .IN1(data_out[18]), .IN2(n70), .IN3(data_in[18]), .IN4(n36), 
        .Q(n50) );
  AO22X1 U23 ( .IN1(data_out[19]), .IN2(n1), .IN3(data_in[19]), .IN4(n36), .Q(
        n49) );
  AO22X1 U24 ( .IN1(data_out[20]), .IN2(n70), .IN3(data_in[20]), .IN4(n36), 
        .Q(n48) );
  AO22X1 U25 ( .IN1(data_out[21]), .IN2(n1), .IN3(data_in[21]), .IN4(n36), .Q(
        n47) );
  AO22X1 U26 ( .IN1(data_out[22]), .IN2(n70), .IN3(data_in[22]), .IN4(n36), 
        .Q(n46) );
  AO22X1 U27 ( .IN1(data_out[23]), .IN2(n1), .IN3(data_in[23]), .IN4(n36), .Q(
        n45) );
  AO22X1 U28 ( .IN1(data_out[24]), .IN2(n70), .IN3(data_in[24]), .IN4(n36), 
        .Q(n44) );
  AO22X1 U29 ( .IN1(data_out[25]), .IN2(n1), .IN3(data_in[25]), .IN4(n36), .Q(
        n43) );
  AO22X1 U30 ( .IN1(data_out[26]), .IN2(n70), .IN3(data_in[26]), .IN4(n36), 
        .Q(n42) );
  AO22X1 U31 ( .IN1(data_out[27]), .IN2(n1), .IN3(data_in[27]), .IN4(n36), .Q(
        n41) );
  AO22X1 U32 ( .IN1(data_out[28]), .IN2(n70), .IN3(data_in[28]), .IN4(n36), 
        .Q(n40) );
  AO22X1 U33 ( .IN1(data_out[29]), .IN2(n1), .IN3(data_in[29]), .IN4(n36), .Q(
        n39) );
  AO22X1 U34 ( .IN1(data_out[30]), .IN2(n70), .IN3(data_in[30]), .IN4(n36), 
        .Q(n38) );
  AO22X1 U35 ( .IN1(data_out[31]), .IN2(n1), .IN3(data_in[31]), .IN4(n36), .Q(
        n37) );
  INVX0 U2 ( .INP(n69), .ZN(n36) );
  AND2X1 U3 ( .IN1(nrst), .IN2(n69), .Q(n70) );
  AND2X1 U36 ( .IN1(nrst), .IN2(n69), .Q(n1) );
  NAND2X1 U37 ( .IN1(nrst), .IN2(en), .QN(n69) );
endmodule


module reg32_2 ( clk, nrst, en, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, nrst, en;
  wire   n1, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71;

  DFFX1 \data_out_reg[31]  ( .D(n38), .CLK(clk), .Q(data_out[31]) );
  DFFX1 \data_out_reg[30]  ( .D(n39), .CLK(clk), .Q(data_out[30]) );
  DFFX1 \data_out_reg[29]  ( .D(n40), .CLK(clk), .Q(data_out[29]) );
  DFFX1 \data_out_reg[28]  ( .D(n41), .CLK(clk), .Q(data_out[28]) );
  DFFX1 \data_out_reg[27]  ( .D(n42), .CLK(clk), .Q(data_out[27]) );
  DFFX1 \data_out_reg[26]  ( .D(n43), .CLK(clk), .Q(data_out[26]) );
  DFFX1 \data_out_reg[25]  ( .D(n44), .CLK(clk), .Q(data_out[25]) );
  DFFX1 \data_out_reg[24]  ( .D(n45), .CLK(clk), .Q(data_out[24]) );
  DFFX1 \data_out_reg[23]  ( .D(n46), .CLK(clk), .Q(data_out[23]) );
  DFFX1 \data_out_reg[22]  ( .D(n47), .CLK(clk), .Q(data_out[22]) );
  DFFX1 \data_out_reg[21]  ( .D(n48), .CLK(clk), .Q(data_out[21]) );
  DFFX1 \data_out_reg[20]  ( .D(n49), .CLK(clk), .Q(data_out[20]) );
  DFFX1 \data_out_reg[19]  ( .D(n50), .CLK(clk), .Q(data_out[19]) );
  DFFX1 \data_out_reg[18]  ( .D(n51), .CLK(clk), .Q(data_out[18]) );
  DFFX1 \data_out_reg[17]  ( .D(n52), .CLK(clk), .Q(data_out[17]) );
  DFFX1 \data_out_reg[16]  ( .D(n53), .CLK(clk), .Q(data_out[16]) );
  DFFX1 \data_out_reg[15]  ( .D(n54), .CLK(clk), .Q(data_out[15]) );
  DFFX1 \data_out_reg[14]  ( .D(n55), .CLK(clk), .Q(data_out[14]) );
  DFFX1 \data_out_reg[13]  ( .D(n56), .CLK(clk), .Q(data_out[13]) );
  DFFX1 \data_out_reg[12]  ( .D(n57), .CLK(clk), .Q(data_out[12]) );
  DFFX1 \data_out_reg[11]  ( .D(n58), .CLK(clk), .Q(data_out[11]) );
  DFFX1 \data_out_reg[10]  ( .D(n59), .CLK(clk), .Q(data_out[10]) );
  DFFX1 \data_out_reg[9]  ( .D(n60), .CLK(clk), .Q(data_out[9]) );
  DFFX1 \data_out_reg[8]  ( .D(n61), .CLK(clk), .Q(data_out[8]) );
  DFFX1 \data_out_reg[7]  ( .D(n62), .CLK(clk), .Q(data_out[7]) );
  DFFX1 \data_out_reg[6]  ( .D(n63), .CLK(clk), .Q(data_out[6]) );
  DFFX1 \data_out_reg[5]  ( .D(n64), .CLK(clk), .Q(data_out[5]) );
  DFFX1 \data_out_reg[4]  ( .D(n65), .CLK(clk), .Q(data_out[4]) );
  DFFX1 \data_out_reg[3]  ( .D(n66), .CLK(clk), .Q(data_out[3]) );
  DFFX1 \data_out_reg[2]  ( .D(n67), .CLK(clk), .Q(data_out[2]) );
  DFFX1 \data_out_reg[1]  ( .D(n68), .CLK(clk), .Q(data_out[1]) );
  DFFX1 \data_out_reg[0]  ( .D(n69), .CLK(clk), .Q(data_out[0]) );
  AO22X1 U4 ( .IN1(data_out[0]), .IN2(n36), .IN3(data_in[0]), .IN4(n37), .Q(
        n69) );
  AO22X1 U5 ( .IN1(data_out[1]), .IN2(n1), .IN3(data_in[1]), .IN4(n37), .Q(n68) );
  AO22X1 U6 ( .IN1(data_out[2]), .IN2(n71), .IN3(data_in[2]), .IN4(n37), .Q(
        n67) );
  AO22X1 U7 ( .IN1(data_out[3]), .IN2(n36), .IN3(data_in[3]), .IN4(n37), .Q(
        n66) );
  AO22X1 U8 ( .IN1(data_out[4]), .IN2(n1), .IN3(data_in[4]), .IN4(n37), .Q(n65) );
  AO22X1 U9 ( .IN1(data_out[5]), .IN2(n71), .IN3(data_in[5]), .IN4(n37), .Q(
        n64) );
  AO22X1 U10 ( .IN1(data_out[6]), .IN2(n36), .IN3(data_in[6]), .IN4(n37), .Q(
        n63) );
  AO22X1 U11 ( .IN1(data_out[7]), .IN2(n1), .IN3(data_in[7]), .IN4(n37), .Q(
        n62) );
  AO22X1 U12 ( .IN1(data_out[8]), .IN2(n71), .IN3(data_in[8]), .IN4(n37), .Q(
        n61) );
  AO22X1 U13 ( .IN1(data_out[9]), .IN2(n36), .IN3(data_in[9]), .IN4(n37), .Q(
        n60) );
  AO22X1 U14 ( .IN1(data_out[10]), .IN2(n1), .IN3(data_in[10]), .IN4(n37), .Q(
        n59) );
  AO22X1 U15 ( .IN1(data_out[11]), .IN2(n71), .IN3(data_in[11]), .IN4(n37), 
        .Q(n58) );
  AO22X1 U16 ( .IN1(data_out[12]), .IN2(n36), .IN3(data_in[12]), .IN4(n37), 
        .Q(n57) );
  AO22X1 U17 ( .IN1(data_out[13]), .IN2(n1), .IN3(data_in[13]), .IN4(n37), .Q(
        n56) );
  AO22X1 U18 ( .IN1(data_out[14]), .IN2(n71), .IN3(data_in[14]), .IN4(n37), 
        .Q(n55) );
  AO22X1 U19 ( .IN1(data_out[15]), .IN2(n36), .IN3(data_in[15]), .IN4(n37), 
        .Q(n54) );
  AO22X1 U20 ( .IN1(data_out[16]), .IN2(n1), .IN3(data_in[16]), .IN4(n37), .Q(
        n53) );
  AO22X1 U21 ( .IN1(data_out[17]), .IN2(n71), .IN3(data_in[17]), .IN4(n37), 
        .Q(n52) );
  AO22X1 U22 ( .IN1(data_out[18]), .IN2(n36), .IN3(data_in[18]), .IN4(n37), 
        .Q(n51) );
  AO22X1 U23 ( .IN1(data_out[19]), .IN2(n1), .IN3(data_in[19]), .IN4(n37), .Q(
        n50) );
  AO22X1 U24 ( .IN1(data_out[20]), .IN2(n71), .IN3(data_in[20]), .IN4(n37), 
        .Q(n49) );
  AO22X1 U25 ( .IN1(data_out[21]), .IN2(n36), .IN3(data_in[21]), .IN4(n37), 
        .Q(n48) );
  AO22X1 U26 ( .IN1(data_out[22]), .IN2(n1), .IN3(data_in[22]), .IN4(n37), .Q(
        n47) );
  AO22X1 U27 ( .IN1(data_out[23]), .IN2(n71), .IN3(data_in[23]), .IN4(n37), 
        .Q(n46) );
  AO22X1 U28 ( .IN1(data_out[24]), .IN2(n36), .IN3(data_in[24]), .IN4(n37), 
        .Q(n45) );
  AO22X1 U29 ( .IN1(data_out[25]), .IN2(n1), .IN3(data_in[25]), .IN4(n37), .Q(
        n44) );
  AO22X1 U30 ( .IN1(data_out[26]), .IN2(n71), .IN3(data_in[26]), .IN4(n37), 
        .Q(n43) );
  AO22X1 U31 ( .IN1(data_out[27]), .IN2(n36), .IN3(data_in[27]), .IN4(n37), 
        .Q(n42) );
  AO22X1 U32 ( .IN1(data_out[28]), .IN2(n1), .IN3(data_in[28]), .IN4(n37), .Q(
        n41) );
  AO22X1 U33 ( .IN1(data_out[29]), .IN2(n71), .IN3(data_in[29]), .IN4(n37), 
        .Q(n40) );
  AO22X1 U34 ( .IN1(data_out[30]), .IN2(n36), .IN3(data_in[30]), .IN4(n37), 
        .Q(n39) );
  AO22X1 U35 ( .IN1(data_out[31]), .IN2(n1), .IN3(data_in[31]), .IN4(n37), .Q(
        n38) );
  INVX0 U2 ( .INP(n70), .ZN(n37) );
  AND2X1 U3 ( .IN1(nrst), .IN2(n70), .Q(n36) );
  AND2X1 U36 ( .IN1(nrst), .IN2(n70), .Q(n1) );
  AND2X1 U37 ( .IN1(nrst), .IN2(n70), .Q(n71) );
  NAND2X1 U38 ( .IN1(nrst), .IN2(en), .QN(n70) );
endmodule


module reg32_1 ( clk, nrst, en, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, nrst, en;
  wire   n1, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71;

  DFFX1 \data_out_reg[31]  ( .D(n38), .CLK(clk), .Q(data_out[31]) );
  DFFX1 \data_out_reg[30]  ( .D(n39), .CLK(clk), .Q(data_out[30]) );
  DFFX1 \data_out_reg[29]  ( .D(n40), .CLK(clk), .Q(data_out[29]) );
  DFFX1 \data_out_reg[28]  ( .D(n41), .CLK(clk), .Q(data_out[28]) );
  DFFX1 \data_out_reg[27]  ( .D(n42), .CLK(clk), .Q(data_out[27]) );
  DFFX1 \data_out_reg[26]  ( .D(n43), .CLK(clk), .Q(data_out[26]) );
  DFFX1 \data_out_reg[25]  ( .D(n44), .CLK(clk), .Q(data_out[25]) );
  DFFX1 \data_out_reg[24]  ( .D(n45), .CLK(clk), .Q(data_out[24]) );
  DFFX1 \data_out_reg[23]  ( .D(n46), .CLK(clk), .Q(data_out[23]) );
  DFFX1 \data_out_reg[22]  ( .D(n47), .CLK(clk), .Q(data_out[22]) );
  DFFX1 \data_out_reg[21]  ( .D(n48), .CLK(clk), .Q(data_out[21]) );
  DFFX1 \data_out_reg[20]  ( .D(n49), .CLK(clk), .Q(data_out[20]) );
  DFFX1 \data_out_reg[19]  ( .D(n50), .CLK(clk), .Q(data_out[19]) );
  DFFX1 \data_out_reg[18]  ( .D(n51), .CLK(clk), .Q(data_out[18]) );
  DFFX1 \data_out_reg[17]  ( .D(n52), .CLK(clk), .Q(data_out[17]) );
  DFFX1 \data_out_reg[16]  ( .D(n53), .CLK(clk), .Q(data_out[16]) );
  DFFX1 \data_out_reg[15]  ( .D(n54), .CLK(clk), .Q(data_out[15]) );
  DFFX1 \data_out_reg[14]  ( .D(n55), .CLK(clk), .Q(data_out[14]) );
  DFFX1 \data_out_reg[13]  ( .D(n56), .CLK(clk), .Q(data_out[13]) );
  DFFX1 \data_out_reg[12]  ( .D(n57), .CLK(clk), .Q(data_out[12]) );
  DFFX1 \data_out_reg[11]  ( .D(n58), .CLK(clk), .Q(data_out[11]) );
  DFFX1 \data_out_reg[10]  ( .D(n59), .CLK(clk), .Q(data_out[10]) );
  DFFX1 \data_out_reg[9]  ( .D(n60), .CLK(clk), .Q(data_out[9]) );
  DFFX1 \data_out_reg[8]  ( .D(n61), .CLK(clk), .Q(data_out[8]) );
  DFFX1 \data_out_reg[7]  ( .D(n62), .CLK(clk), .Q(data_out[7]) );
  DFFX1 \data_out_reg[6]  ( .D(n63), .CLK(clk), .Q(data_out[6]) );
  DFFX1 \data_out_reg[5]  ( .D(n64), .CLK(clk), .Q(data_out[5]) );
  DFFX1 \data_out_reg[4]  ( .D(n65), .CLK(clk), .Q(data_out[4]) );
  DFFX1 \data_out_reg[3]  ( .D(n66), .CLK(clk), .Q(data_out[3]) );
  DFFX1 \data_out_reg[2]  ( .D(n67), .CLK(clk), .Q(data_out[2]) );
  DFFX1 \data_out_reg[1]  ( .D(n68), .CLK(clk), .Q(data_out[1]) );
  DFFX1 \data_out_reg[0]  ( .D(n69), .CLK(clk), .Q(data_out[0]) );
  AO22X1 U4 ( .IN1(data_out[0]), .IN2(n36), .IN3(data_in[0]), .IN4(n37), .Q(
        n69) );
  AO22X1 U5 ( .IN1(data_out[1]), .IN2(n1), .IN3(data_in[1]), .IN4(n37), .Q(n68) );
  AO22X1 U6 ( .IN1(data_out[2]), .IN2(n71), .IN3(data_in[2]), .IN4(n37), .Q(
        n67) );
  AO22X1 U7 ( .IN1(data_out[3]), .IN2(n36), .IN3(data_in[3]), .IN4(n37), .Q(
        n66) );
  AO22X1 U8 ( .IN1(data_out[4]), .IN2(n1), .IN3(data_in[4]), .IN4(n37), .Q(n65) );
  AO22X1 U9 ( .IN1(data_out[5]), .IN2(n71), .IN3(data_in[5]), .IN4(n37), .Q(
        n64) );
  AO22X1 U10 ( .IN1(data_out[6]), .IN2(n36), .IN3(data_in[6]), .IN4(n37), .Q(
        n63) );
  AO22X1 U11 ( .IN1(data_out[7]), .IN2(n1), .IN3(data_in[7]), .IN4(n37), .Q(
        n62) );
  AO22X1 U12 ( .IN1(data_out[8]), .IN2(n71), .IN3(data_in[8]), .IN4(n37), .Q(
        n61) );
  AO22X1 U13 ( .IN1(data_out[9]), .IN2(n36), .IN3(data_in[9]), .IN4(n37), .Q(
        n60) );
  AO22X1 U14 ( .IN1(data_out[10]), .IN2(n1), .IN3(data_in[10]), .IN4(n37), .Q(
        n59) );
  AO22X1 U15 ( .IN1(data_out[11]), .IN2(n71), .IN3(data_in[11]), .IN4(n37), 
        .Q(n58) );
  AO22X1 U16 ( .IN1(data_out[12]), .IN2(n36), .IN3(data_in[12]), .IN4(n37), 
        .Q(n57) );
  AO22X1 U17 ( .IN1(data_out[13]), .IN2(n1), .IN3(data_in[13]), .IN4(n37), .Q(
        n56) );
  AO22X1 U18 ( .IN1(data_out[14]), .IN2(n71), .IN3(data_in[14]), .IN4(n37), 
        .Q(n55) );
  AO22X1 U19 ( .IN1(data_out[15]), .IN2(n36), .IN3(data_in[15]), .IN4(n37), 
        .Q(n54) );
  AO22X1 U20 ( .IN1(data_out[16]), .IN2(n1), .IN3(data_in[16]), .IN4(n37), .Q(
        n53) );
  AO22X1 U21 ( .IN1(data_out[17]), .IN2(n71), .IN3(data_in[17]), .IN4(n37), 
        .Q(n52) );
  AO22X1 U22 ( .IN1(data_out[18]), .IN2(n36), .IN3(data_in[18]), .IN4(n37), 
        .Q(n51) );
  AO22X1 U23 ( .IN1(data_out[19]), .IN2(n1), .IN3(data_in[19]), .IN4(n37), .Q(
        n50) );
  AO22X1 U24 ( .IN1(data_out[20]), .IN2(n71), .IN3(data_in[20]), .IN4(n37), 
        .Q(n49) );
  AO22X1 U25 ( .IN1(data_out[21]), .IN2(n36), .IN3(data_in[21]), .IN4(n37), 
        .Q(n48) );
  AO22X1 U26 ( .IN1(data_out[22]), .IN2(n1), .IN3(data_in[22]), .IN4(n37), .Q(
        n47) );
  AO22X1 U27 ( .IN1(data_out[23]), .IN2(n71), .IN3(data_in[23]), .IN4(n37), 
        .Q(n46) );
  AO22X1 U28 ( .IN1(data_out[24]), .IN2(n36), .IN3(data_in[24]), .IN4(n37), 
        .Q(n45) );
  AO22X1 U29 ( .IN1(data_out[25]), .IN2(n1), .IN3(data_in[25]), .IN4(n37), .Q(
        n44) );
  AO22X1 U30 ( .IN1(data_out[26]), .IN2(n71), .IN3(data_in[26]), .IN4(n37), 
        .Q(n43) );
  AO22X1 U31 ( .IN1(data_out[27]), .IN2(n36), .IN3(data_in[27]), .IN4(n37), 
        .Q(n42) );
  AO22X1 U32 ( .IN1(data_out[28]), .IN2(n1), .IN3(data_in[28]), .IN4(n37), .Q(
        n41) );
  AO22X1 U33 ( .IN1(data_out[29]), .IN2(n71), .IN3(data_in[29]), .IN4(n37), 
        .Q(n40) );
  AO22X1 U34 ( .IN1(data_out[30]), .IN2(n36), .IN3(data_in[30]), .IN4(n37), 
        .Q(n39) );
  AO22X1 U35 ( .IN1(data_out[31]), .IN2(n1), .IN3(data_in[31]), .IN4(n37), .Q(
        n38) );
  INVX0 U2 ( .INP(n70), .ZN(n37) );
  AND2X1 U3 ( .IN1(nrst), .IN2(n70), .Q(n36) );
  AND2X1 U36 ( .IN1(nrst), .IN2(n70), .Q(n1) );
  AND2X1 U37 ( .IN1(nrst), .IN2(n70), .Q(n71) );
  NAND2X1 U38 ( .IN1(nrst), .IN2(en), .QN(n70) );
endmodule


module control ( clk, nrst, zero, inst, jr, jal, jal_pc, load, wr_mem, use_imm, 
        sw, debug_inst, alu_code, sel_pc, flush, wr_rf, stall, fwd_opA, 
        fwd_opB, fwd_sw, fwd_jr );
  input [31:0] inst;
  output [159:0] debug_inst;
  output [6:0] alu_code;
  output [2:0] sel_pc;
  output [1:0] flush;
  output [2:0] fwd_opA;
  output [2:0] fwd_opB;
  output [2:0] fwd_sw;
  output [2:0] fwd_jr;
  input clk, nrst, zero;
  output jr, jal, jal_pc, load, wr_mem, use_imm, sw, wr_rf, stall;
  wire   \inst[31] , \inst[30] , \inst[29] , \inst[28] , \inst[27] ,
         \inst[26] , \inst[25] , \inst[24] , \inst[23] , \inst[22] ,
         \inst[21] , \inst[20] , \inst[19] , \inst[18] , \inst[17] ,
         \inst[16] , \inst[15] , \inst[14] , \inst[13] , \inst[12] ,
         \inst[11] , \inst[10] , \inst[9] , \inst[8] , \inst[7] , \inst[6] ,
         \inst[5] , \inst[4] , \inst[3] , \inst[2] , \inst[1] , \inst[0] , jr,
         _5_net_, _7_net_, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n43, n44, n45, n46, n47, n181;
  assign debug_inst[31] = \inst[31] ;
  assign \inst[31]  = inst[31];
  assign debug_inst[30] = \inst[30] ;
  assign \inst[30]  = inst[30];
  assign debug_inst[29] = \inst[29] ;
  assign \inst[29]  = inst[29];
  assign debug_inst[28] = \inst[28] ;
  assign \inst[28]  = inst[28];
  assign debug_inst[27] = \inst[27] ;
  assign \inst[27]  = inst[27];
  assign debug_inst[26] = \inst[26] ;
  assign \inst[26]  = inst[26];
  assign debug_inst[25] = \inst[25] ;
  assign \inst[25]  = inst[25];
  assign debug_inst[24] = \inst[24] ;
  assign \inst[24]  = inst[24];
  assign debug_inst[23] = \inst[23] ;
  assign \inst[23]  = inst[23];
  assign debug_inst[22] = \inst[22] ;
  assign \inst[22]  = inst[22];
  assign debug_inst[21] = \inst[21] ;
  assign \inst[21]  = inst[21];
  assign debug_inst[20] = \inst[20] ;
  assign \inst[20]  = inst[20];
  assign debug_inst[19] = \inst[19] ;
  assign \inst[19]  = inst[19];
  assign debug_inst[18] = \inst[18] ;
  assign \inst[18]  = inst[18];
  assign debug_inst[17] = \inst[17] ;
  assign \inst[17]  = inst[17];
  assign debug_inst[16] = \inst[16] ;
  assign \inst[16]  = inst[16];
  assign debug_inst[15] = \inst[15] ;
  assign \inst[15]  = inst[15];
  assign debug_inst[14] = \inst[14] ;
  assign \inst[14]  = inst[14];
  assign debug_inst[13] = \inst[13] ;
  assign \inst[13]  = inst[13];
  assign debug_inst[12] = \inst[12] ;
  assign \inst[12]  = inst[12];
  assign debug_inst[11] = \inst[11] ;
  assign \inst[11]  = inst[11];
  assign debug_inst[10] = \inst[10] ;
  assign \inst[10]  = inst[10];
  assign debug_inst[9] = \inst[9] ;
  assign \inst[9]  = inst[9];
  assign debug_inst[8] = \inst[8] ;
  assign \inst[8]  = inst[8];
  assign debug_inst[7] = \inst[7] ;
  assign \inst[7]  = inst[7];
  assign debug_inst[6] = \inst[6] ;
  assign \inst[6]  = inst[6];
  assign debug_inst[5] = \inst[5] ;
  assign \inst[5]  = inst[5];
  assign debug_inst[4] = \inst[4] ;
  assign \inst[4]  = inst[4];
  assign debug_inst[3] = \inst[3] ;
  assign \inst[3]  = inst[3];
  assign debug_inst[2] = \inst[2] ;
  assign \inst[2]  = inst[2];
  assign debug_inst[1] = \inst[1] ;
  assign \inst[1]  = inst[1];
  assign debug_inst[0] = \inst[0] ;
  assign \inst[0]  = inst[0];
  assign sel_pc[0] = jr;

  OR3X1 U94 ( .IN1(n50), .IN2(n51), .IN3(n47), .Q(n49) );
  NOR3X0 U95 ( .IN1(debug_inst[34]), .IN2(debug_inst[36]), .IN3(n52), .QN(
        use_imm) );
  AND2X1 U96 ( .IN1(n53), .IN2(n54), .Q(n52) );
  OR3X1 U97 ( .IN1(debug_inst[32]), .IN2(debug_inst[37]), .IN3(n26), .Q(n54)
         );
  AND2X1 U98 ( .IN1(n30), .IN2(debug_inst[95]), .Q(alu_code[6]) );
  OA221X1 U99 ( .IN1(n68), .IN2(n39), .IN3(n69), .IN4(n36), .IN5(n70), .Q(n67)
         );
  AND2X1 U100 ( .IN1(n30), .IN2(debug_inst[93]), .Q(alu_code[4]) );
  AO22X1 U101 ( .IN1(n75), .IN2(n38), .IN3(n30), .IN4(debug_inst[92]), .Q(
        alu_code[3]) );
  AND2X1 U102 ( .IN1(n30), .IN2(debug_inst[91]), .Q(alu_code[2]) );
  OAI22X1 U103 ( .IN1(n31), .IN2(n76), .IN3(n72), .IN4(debug_inst[68]), .QN(
        alu_code[1]) );
  NOR3X0 U104 ( .IN1(n78), .IN2(debug_inst[64]), .IN3(n39), .QN(n75) );
  NOR3X0 U105 ( .IN1(n3), .IN2(stall), .IN3(sel_pc[2]), .QN(_7_net_) );
  AO21X1 U106 ( .IN1(n79), .IN2(n5), .IN3(flush[0]), .Q(flush[1]) );
  AND2X1 U107 ( .IN1(sel_pc[2]), .IN2(n5), .Q(flush[0]) );
  AND3X1 U108 ( .IN1(n80), .IN2(n38), .IN3(n77), .Q(sel_pc[2]) );
  NOR4X0 U109 ( .IN1(n40), .IN2(debug_inst[65]), .IN3(debug_inst[67]), .IN4(
        debug_inst[69]), .QN(n77) );
  XOR2X1 U110 ( .IN1(zero), .IN2(debug_inst[64]), .Q(n80) );
  AO222X1 U111 ( .IN1(debug_inst[133]), .IN2(n81), .IN3(n37), .IN4(n82), .IN5(
        load), .IN6(n83), .Q(stall) );
  NAND3X0 U112 ( .IN1(n60), .IN2(n57), .IN3(n63), .QN(n83) );
  NAND4X0 U113 ( .IN1(n84), .IN2(n85), .IN3(n86), .IN4(n87), .QN(n63) );
  NOR4X0 U114 ( .IN1(n88), .IN2(n89), .IN3(n90), .IN4(n91), .QN(n87) );
  XOR2X1 U115 ( .IN1(n21), .IN2(n92), .Q(n91) );
  XNOR2X1 U116 ( .IN1(debug_inst[38]), .IN2(n93), .Q(n89) );
  XOR2X1 U117 ( .IN1(n94), .IN2(debug_inst[39]), .Q(n86) );
  XOR2X1 U118 ( .IN1(n95), .IN2(debug_inst[41]), .Q(n85) );
  XOR2X1 U119 ( .IN1(n96), .IN2(debug_inst[40]), .Q(n84) );
  NAND4X0 U120 ( .IN1(n97), .IN2(n98), .IN3(n99), .IN4(n100), .QN(n57) );
  NOR4X0 U121 ( .IN1(n88), .IN2(n101), .IN3(n102), .IN4(n103), .QN(n100) );
  XOR2X1 U122 ( .IN1(n15), .IN2(n92), .Q(n103) );
  XNOR2X1 U123 ( .IN1(debug_inst[52]), .IN2(n93), .Q(n101) );
  XOR2X1 U124 ( .IN1(n94), .IN2(debug_inst[53]), .Q(n99) );
  XOR2X1 U125 ( .IN1(n95), .IN2(debug_inst[55]), .Q(n98) );
  XOR2X1 U126 ( .IN1(n96), .IN2(debug_inst[54]), .Q(n97) );
  NAND4X0 U127 ( .IN1(n104), .IN2(n105), .IN3(n106), .IN4(n107), .QN(n60) );
  NOR4X0 U128 ( .IN1(n88), .IN2(n108), .IN3(n109), .IN4(n110), .QN(n107) );
  XOR2X1 U129 ( .IN1(n18), .IN2(n92), .Q(n110) );
  XNOR2X1 U130 ( .IN1(debug_inst[47]), .IN2(n93), .Q(n108) );
  NOR3X0 U131 ( .IN1(jal_pc), .IN2(load), .IN3(n112), .QN(n88) );
  AND4X1 U132 ( .IN1(n113), .IN2(n43), .IN3(n114), .IN4(n41), .Q(n112) );
  AO21X1 U133 ( .IN1(n115), .IN2(n45), .IN3(debug_inst[99]), .Q(n113) );
  NAND3X0 U134 ( .IN1(n116), .IN2(debug_inst[124]), .IN3(n117), .QN(n115) );
  NOR4X0 U135 ( .IN1(debug_inst[127]), .IN2(debug_inst[126]), .IN3(
        debug_inst[125]), .IN4(debug_inst[123]), .QN(n117) );
  XOR2X1 U136 ( .IN1(n94), .IN2(debug_inst[48]), .Q(n106) );
  XOR2X1 U137 ( .IN1(n95), .IN2(debug_inst[50]), .Q(n105) );
  XOR2X1 U138 ( .IN1(n96), .IN2(debug_inst[49]), .Q(n104) );
  NAND4X0 U139 ( .IN1(debug_inst[96]), .IN2(n43), .IN3(debug_inst[97]), .IN4(
        n118), .QN(n111) );
  NOR3X0 U140 ( .IN1(debug_inst[101]), .IN2(debug_inst[99]), .IN3(
        debug_inst[98]), .QN(n118) );
  NAND4X0 U141 ( .IN1(debug_inst[97]), .IN2(debug_inst[96]), .IN3(n119), .IN4(
        debug_inst[101]), .QN(n65) );
  NAND3X0 U142 ( .IN1(n59), .IN2(n56), .IN3(n62), .QN(n82) );
  NAND4X0 U143 ( .IN1(n120), .IN2(n121), .IN3(n122), .IN4(n123), .QN(n62) );
  NOR4X0 U144 ( .IN1(n124), .IN2(n125), .IN3(n90), .IN4(n126), .QN(n123) );
  XOR2X1 U145 ( .IN1(n21), .IN2(n127), .Q(n126) );
  XNOR2X1 U146 ( .IN1(debug_inst[38]), .IN2(n128), .Q(n125) );
  XOR2X1 U147 ( .IN1(n129), .IN2(debug_inst[39]), .Q(n122) );
  XOR2X1 U148 ( .IN1(n130), .IN2(debug_inst[41]), .Q(n121) );
  XOR2X1 U149 ( .IN1(n131), .IN2(debug_inst[40]), .Q(n120) );
  NAND4X0 U150 ( .IN1(n132), .IN2(n133), .IN3(n134), .IN4(n135), .QN(n56) );
  NOR4X0 U151 ( .IN1(n124), .IN2(n136), .IN3(n102), .IN4(n137), .QN(n135) );
  XOR2X1 U152 ( .IN1(n15), .IN2(n127), .Q(n137) );
  XNOR2X1 U153 ( .IN1(debug_inst[52]), .IN2(n128), .Q(n136) );
  XOR2X1 U154 ( .IN1(n129), .IN2(debug_inst[53]), .Q(n134) );
  XOR2X1 U155 ( .IN1(n130), .IN2(debug_inst[55]), .Q(n133) );
  XOR2X1 U156 ( .IN1(n131), .IN2(debug_inst[54]), .Q(n132) );
  NAND4X0 U157 ( .IN1(n138), .IN2(n139), .IN3(n140), .IN4(n141), .QN(n59) );
  NOR4X0 U158 ( .IN1(n124), .IN2(n142), .IN3(n109), .IN4(n143), .QN(n141) );
  XOR2X1 U159 ( .IN1(n18), .IN2(n127), .Q(n143) );
  XNOR2X1 U160 ( .IN1(debug_inst[47]), .IN2(n128), .Q(n142) );
  AND3X1 U161 ( .IN1(n144), .IN2(n76), .IN3(n145), .Q(n124) );
  NAND3X0 U162 ( .IN1(n40), .IN2(n38), .IN3(n146), .QN(n145) );
  AO22X1 U163 ( .IN1(n37), .IN2(n39), .IN3(n147), .IN4(debug_inst[67]), .Q(
        n146) );
  NAND3X0 U164 ( .IN1(n74), .IN2(n38), .IN3(n73), .QN(n76) );
  OR4X1 U165 ( .IN1(debug_inst[64]), .IN2(debug_inst[65]), .IN3(debug_inst[66]), .IN4(debug_inst[69]), .Q(n68) );
  NAND4X0 U166 ( .IN1(n32), .IN2(n31), .IN3(debug_inst[92]), .IN4(n148), .QN(
        n74) );
  NOR4X0 U167 ( .IN1(debug_inst[95]), .IN2(debug_inst[94]), .IN3(
        debug_inst[93]), .IN4(debug_inst[91]), .QN(n148) );
  XOR2X1 U168 ( .IN1(n129), .IN2(debug_inst[48]), .Q(n140) );
  XOR2X1 U169 ( .IN1(n130), .IN2(debug_inst[50]), .Q(n139) );
  XOR2X1 U170 ( .IN1(n131), .IN2(debug_inst[49]), .Q(n138) );
  NAND4X0 U171 ( .IN1(n34), .IN2(debug_inst[64]), .IN3(n39), .IN4(n38), .QN(
        n144) );
  NAND3X0 U172 ( .IN1(n40), .IN2(n35), .IN3(debug_inst[65]), .QN(n78) );
  NAND3X0 U173 ( .IN1(debug_inst[65]), .IN2(debug_inst[64]), .IN3(
        debug_inst[69]), .QN(n71) );
  NAND3X0 U174 ( .IN1(n61), .IN2(n58), .IN3(n64), .QN(n81) );
  NAND4X0 U175 ( .IN1(n149), .IN2(n150), .IN3(n151), .IN4(n152), .QN(n64) );
  NOR4X0 U176 ( .IN1(n153), .IN2(n154), .IN3(n90), .IN4(n155), .QN(n152) );
  XOR2X1 U177 ( .IN1(n21), .IN2(n156), .Q(n155) );
  NAND4X0 U178 ( .IN1(n22), .IN2(n21), .IN3(n23), .IN4(n159), .QN(n158) );
  AO21X1 U179 ( .IN1(n11), .IN2(n79), .IN3(sw), .Q(n157) );
  NOR4X0 U180 ( .IN1(n53), .IN2(n26), .IN3(debug_inst[34]), .IN4(
        debug_inst[36]), .QN(sw) );
  NAND3X0 U181 ( .IN1(debug_inst[33]), .IN2(debug_inst[32]), .IN3(
        debug_inst[37]), .QN(n53) );
  XOR2X1 U182 ( .IN1(n160), .IN2(debug_inst[38]), .Q(n154) );
  XOR2X1 U183 ( .IN1(n161), .IN2(debug_inst[39]), .Q(n151) );
  XOR2X1 U184 ( .IN1(n162), .IN2(debug_inst[41]), .Q(n150) );
  XOR2X1 U185 ( .IN1(n163), .IN2(debug_inst[40]), .Q(n149) );
  NAND4X0 U186 ( .IN1(n164), .IN2(n165), .IN3(n166), .IN4(n167), .QN(n58) );
  NOR4X0 U187 ( .IN1(n153), .IN2(n168), .IN3(n102), .IN4(n169), .QN(n167) );
  XOR2X1 U188 ( .IN1(n15), .IN2(n156), .Q(n169) );
  NAND4X0 U189 ( .IN1(n170), .IN2(n171), .IN3(n172), .IN4(n27), .QN(n102) );
  AO21X1 U190 ( .IN1(n173), .IN2(n28), .IN3(debug_inst[34]), .Q(n172) );
  NAND4X0 U191 ( .IN1(n16), .IN2(n15), .IN3(n17), .IN4(n174), .QN(n171) );
  XOR2X1 U192 ( .IN1(n160), .IN2(debug_inst[52]), .Q(n168) );
  XOR2X1 U193 ( .IN1(n161), .IN2(debug_inst[53]), .Q(n166) );
  XOR2X1 U194 ( .IN1(n162), .IN2(debug_inst[55]), .Q(n165) );
  XOR2X1 U195 ( .IN1(n163), .IN2(debug_inst[54]), .Q(n164) );
  NAND4X0 U196 ( .IN1(n175), .IN2(n176), .IN3(n177), .IN4(n178), .QN(n61) );
  NOR4X0 U197 ( .IN1(n153), .IN2(n179), .IN3(n109), .IN4(n180), .QN(n178) );
  XOR2X1 U198 ( .IN1(n18), .IN2(n156), .Q(n180) );
  XOR2X1 U200 ( .IN1(n160), .IN2(debug_inst[47]), .Q(n179) );
  OR2X1 U201 ( .IN1(n183), .IN2(debug_inst[134]), .Q(n160) );
  OR2X1 U202 ( .IN1(debug_inst[128]), .IN2(debug_inst[133]), .Q(n50) );
  OR4X1 U203 ( .IN1(n186), .IN2(debug_inst[129]), .IN3(debug_inst[130]), .IN4(
        debug_inst[132]), .Q(n185) );
  AND3X1 U204 ( .IN1(n187), .IN2(debug_inst[156]), .IN3(n188), .Q(n186) );
  NOR4X0 U205 ( .IN1(debug_inst[159]), .IN2(debug_inst[158]), .IN3(
        debug_inst[157]), .IN4(debug_inst[155]), .QN(n188) );
  XOR2X1 U206 ( .IN1(n161), .IN2(debug_inst[48]), .Q(n177) );
  XOR2X1 U207 ( .IN1(n162), .IN2(debug_inst[50]), .Q(n176) );
  XOR2X1 U208 ( .IN1(n163), .IN2(debug_inst[49]), .Q(n175) );
  NAND3X0 U209 ( .IN1(n51), .IN2(n189), .IN3(debug_inst[128]), .QN(n48) );
  AND2X1 U210 ( .IN1(debug_inst[129]), .IN2(n181), .Q(n51) );
  NAND3X0 U211 ( .IN1(n11), .IN2(n28), .IN3(n190), .QN(n66) );
  NAND3X0 U212 ( .IN1(n191), .IN2(debug_inst[60]), .IN3(n192), .QN(n173) );
  NOR4X0 U213 ( .IN1(debug_inst[63]), .IN2(debug_inst[62]), .IN3(
        debug_inst[61]), .IN4(debug_inst[59]), .QN(n192) );
  NOR3X0 U214 ( .IN1(debug_inst[36]), .IN2(debug_inst[37]), .IN3(
        debug_inst[35]), .QN(n170) );
  reg_fwd FWD_VECTOR ( .clk(clk), .nrst(n2), .fwd_opA0({n6, n7, n4}), 
        .fwd_opB0({n13, n14, n12}), .fwd_jr0({n9, n10, n8}), .fwd_opA(fwd_opA), 
        .fwd_opB(fwd_opB), .fwd_sw(fwd_sw), .fwd_jr(fwd_jr) );
  reg32_4 if_id ( .clk(clk), .nrst(_5_net_), .en(n5), .data_in({\inst[31] , 
        \inst[30] , \inst[29] , \inst[28] , \inst[27] , \inst[26] , \inst[25] , 
        \inst[24] , \inst[23] , \inst[22] , \inst[21] , \inst[20] , \inst[19] , 
        \inst[18] , \inst[17] , \inst[16] , \inst[15] , \inst[14] , \inst[13] , 
        \inst[12] , \inst[11] , \inst[10] , \inst[9] , \inst[8] , \inst[7] , 
        \inst[6] , \inst[5] , \inst[4] , \inst[3] , \inst[2] , \inst[1] , 
        \inst[0] }), .data_out(debug_inst[63:32]) );
  reg32_3 id_exe ( .clk(clk), .nrst(_7_net_), .en(1'b1), .data_in(
        debug_inst[63:32]), .data_out(debug_inst[95:64]) );
  reg32_2 exe_mem ( .clk(clk), .nrst(n2), .en(1'b1), .data_in(
        debug_inst[95:64]), .data_out(debug_inst[127:96]) );
  reg32_1 mem_wb ( .clk(clk), .nrst(n2), .en(1'b1), .data_in(
        debug_inst[127:96]), .data_out(debug_inst[159:128]) );
  INVX0 U3 ( .INP(debug_inst[50]), .ZN(n19) );
  INVX0 U4 ( .INP(n76), .ZN(n30) );
  INVX0 U5 ( .INP(n3), .ZN(n2) );
  NOR2X0 U6 ( .IN1(flush[1]), .IN2(n3), .QN(_5_net_) );
  INVX0 U7 ( .INP(n61), .ZN(n4) );
  INVX0 U8 ( .INP(n60), .ZN(n7) );
  INVX0 U9 ( .INP(n59), .ZN(n6) );
  INVX0 U10 ( .INP(n58), .ZN(n12) );
  INVX0 U11 ( .INP(n57), .ZN(n14) );
  INVX0 U12 ( .INP(n56), .ZN(n13) );
  NOR2X0 U13 ( .IN1(n77), .IN2(n75), .QN(n72) );
  INVX0 U14 ( .INP(n74), .ZN(n29) );
  INVX0 U15 ( .INP(n111), .ZN(jal_pc) );
  INVX0 U16 ( .INP(n183), .ZN(n46) );
  NOR2X0 U17 ( .IN1(n28), .IN2(n55), .QN(jal) );
  INVX0 U18 ( .INP(n63), .ZN(n10) );
  INVX0 U19 ( .INP(n62), .ZN(n9) );
  INVX0 U20 ( .INP(n64), .ZN(n8) );
  NAND2X1 U21 ( .IN1(n55), .IN2(n66), .QN(n79) );
  INVX0 U22 ( .INP(stall), .ZN(n5) );
  INVX0 U23 ( .INP(n55), .ZN(sel_pc[1]) );
  INVX0 U24 ( .INP(n173), .ZN(n11) );
  INVX0 U25 ( .INP(n71), .ZN(n37) );
  INVX0 U26 ( .INP(n189), .ZN(n47) );
  NOR2X0 U27 ( .IN1(debug_inst[98]), .IN2(debug_inst[100]), .QN(n119) );
  NAND2X1 U28 ( .IN1(n48), .IN2(n49), .QN(wr_rf) );
  NOR2X0 U29 ( .IN1(n65), .IN2(n44), .QN(wr_mem) );
  INVX0 U30 ( .INP(debug_inst[99]), .ZN(n44) );
  INVX0 U31 ( .INP(nrst), .ZN(n3) );
  NOR2X0 U32 ( .IN1(n76), .IN2(n32), .QN(alu_code[0]) );
  INVX0 U33 ( .INP(debug_inst[69]), .ZN(n35) );
  INVX0 U34 ( .INP(debug_inst[68]), .ZN(n38) );
  NOR2X0 U35 ( .IN1(n68), .IN2(debug_inst[67]), .QN(n73) );
  INVX0 U36 ( .INP(debug_inst[67]), .ZN(n39) );
  INVX0 U37 ( .INP(debug_inst[66]), .ZN(n40) );
  NOR2X0 U38 ( .IN1(debug_inst[68]), .IN2(n67), .QN(alu_code[5]) );
  INVX0 U39 ( .INP(n73), .ZN(n36) );
  NOR2X0 U40 ( .IN1(n29), .IN2(debug_inst[94]), .QN(n69) );
  INVX0 U41 ( .INP(debug_inst[89]), .ZN(n32) );
  OA21X1 U42 ( .IN1(debug_inst[66]), .IN2(n71), .IN3(n72), .Q(n70) );
  INVX0 U43 ( .INP(debug_inst[90]), .ZN(n31) );
  NOR2X0 U44 ( .IN1(n65), .IN2(debug_inst[99]), .QN(load) );
  INVX0 U45 ( .INP(n78), .ZN(n34) );
  INVX0 U46 ( .INP(debug_inst[101]), .ZN(n41) );
  NOR2X0 U47 ( .IN1(debug_inst[98]), .IN2(debug_inst[96]), .QN(n114) );
  INVX0 U48 ( .INP(debug_inst[33]), .ZN(n27) );
  NAND2X1 U49 ( .IN1(debug_inst[71]), .IN2(n144), .QN(n129) );
  NAND2X1 U50 ( .IN1(debug_inst[73]), .IN2(n144), .QN(n130) );
  NAND2X1 U51 ( .IN1(debug_inst[72]), .IN2(n144), .QN(n131) );
  NAND2X1 U52 ( .IN1(debug_inst[103]), .IN2(n111), .QN(n94) );
  NAND2X1 U53 ( .IN1(debug_inst[105]), .IN2(n111), .QN(n95) );
  NAND2X1 U54 ( .IN1(debug_inst[104]), .IN2(n111), .QN(n96) );
  NAND2X1 U55 ( .IN1(debug_inst[74]), .IN2(n144), .QN(n127) );
  NAND2X1 U56 ( .IN1(debug_inst[106]), .IN2(n111), .QN(n92) );
  NOR2X0 U57 ( .IN1(debug_inst[58]), .IN2(debug_inst[57]), .QN(n191) );
  NOR2X0 U58 ( .IN1(jal_pc), .IN2(debug_inst[102]), .QN(n93) );
  NOR2X0 U59 ( .IN1(n33), .IN2(debug_inst[70]), .QN(n128) );
  INVX0 U60 ( .INP(n144), .ZN(n33) );
  NOR2X0 U61 ( .IN1(n66), .IN2(debug_inst[33]), .QN(jr) );
  NOR2X0 U62 ( .IN1(debug_inst[69]), .IN2(debug_inst[64]), .QN(n147) );
  NAND2X1 U63 ( .IN1(n190), .IN2(debug_inst[33]), .QN(n55) );
  INVX0 U64 ( .INP(debug_inst[42]), .ZN(n21) );
  INVX0 U65 ( .INP(debug_inst[56]), .ZN(n15) );
  INVX0 U66 ( .INP(debug_inst[51]), .ZN(n18) );
  NOR2X0 U67 ( .IN1(n48), .IN2(debug_inst[133]), .QN(n183) );
  NAND2X1 U68 ( .IN1(debug_inst[135]), .IN2(n46), .QN(n161) );
  NAND2X1 U69 ( .IN1(debug_inst[137]), .IN2(n46), .QN(n162) );
  NAND2X1 U70 ( .IN1(debug_inst[136]), .IN2(n46), .QN(n163) );
  NOR2X0 U71 ( .IN1(n25), .IN2(debug_inst[34]), .QN(n190) );
  INVX0 U72 ( .INP(n170), .ZN(n25) );
  NAND2X1 U73 ( .IN1(debug_inst[138]), .IN2(n46), .QN(n156) );
  NAND2X1 U74 ( .IN1(n157), .IN2(n158), .QN(n90) );
  INVX0 U75 ( .INP(debug_inst[41]), .ZN(n22) );
  OR2X1 U76 ( .IN1(n79), .IN2(n1), .Q(n109) );
  AND4X1 U77 ( .IN1(n19), .IN2(n18), .IN3(n20), .IN4(n182), .Q(n1) );
  INVX0 U78 ( .INP(debug_inst[32]), .ZN(n28) );
  NOR2X0 U79 ( .IN1(debug_inst[39]), .IN2(debug_inst[38]), .QN(n159) );
  NOR2X0 U80 ( .IN1(debug_inst[53]), .IN2(debug_inst[52]), .QN(n174) );
  NOR2X0 U81 ( .IN1(debug_inst[130]), .IN2(debug_inst[132]), .QN(n189) );
  NOR2X0 U82 ( .IN1(debug_inst[48]), .IN2(debug_inst[47]), .QN(n182) );
  OA21X1 U83 ( .IN1(n184), .IN2(n50), .IN3(n48), .Q(n153) );
  OA21X1 U84 ( .IN1(n47), .IN2(n181), .IN3(n185), .Q(n184) );
  INVX0 U85 ( .INP(debug_inst[35]), .ZN(n26) );
  NOR2X0 U86 ( .IN1(debug_inst[154]), .IN2(debug_inst[153]), .QN(n187) );
  INVX0 U87 ( .INP(debug_inst[40]), .ZN(n23) );
  INVX0 U88 ( .INP(debug_inst[97]), .ZN(n45) );
  NOR2X0 U89 ( .IN1(debug_inst[122]), .IN2(debug_inst[121]), .QN(n116) );
  INVX0 U90 ( .INP(debug_inst[54]), .ZN(n17) );
  INVX0 U91 ( .INP(debug_inst[55]), .ZN(n16) );
  INVX0 U92 ( .INP(debug_inst[49]), .ZN(n20) );
  INVX0 U93 ( .INP(debug_inst[100]), .ZN(n43) );
  INVX0 U199 ( .INP(debug_inst[131]), .ZN(n181) );
endmodule


module pipeline_riscv_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(B[0]), .IN2(A[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module pipeline_riscv_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2X1 U1 ( .IN1(A[2]), .IN2(A[3]), .Q(n1) );
  AND2X1 U2 ( .IN1(n1), .IN2(A[4]), .Q(n2) );
  AND2X1 U3 ( .IN1(n2), .IN2(A[5]), .Q(n3) );
  AND2X1 U4 ( .IN1(n3), .IN2(A[6]), .Q(n4) );
  AND2X1 U5 ( .IN1(n4), .IN2(A[7]), .Q(n5) );
  AND2X1 U6 ( .IN1(n5), .IN2(A[8]), .Q(n6) );
  AND2X1 U7 ( .IN1(n6), .IN2(A[9]), .Q(n7) );
  AND2X1 U8 ( .IN1(n7), .IN2(A[10]), .Q(n8) );
  AND2X1 U9 ( .IN1(n8), .IN2(A[11]), .Q(n9) );
  AND2X1 U10 ( .IN1(n9), .IN2(A[12]), .Q(n10) );
  AND2X1 U11 ( .IN1(n10), .IN2(A[13]), .Q(n11) );
  AND2X1 U12 ( .IN1(n11), .IN2(A[14]), .Q(n12) );
  AND2X1 U13 ( .IN1(n12), .IN2(A[15]), .Q(n13) );
  XNOR2X1 U14 ( .IN1(n28), .IN2(A[31]), .Q(SUM[31]) );
  NAND2X1 U15 ( .IN1(n27), .IN2(A[30]), .QN(n28) );
  AND2X1 U16 ( .IN1(n13), .IN2(A[16]), .Q(n14) );
  AND2X1 U17 ( .IN1(n14), .IN2(A[17]), .Q(n15) );
  AND2X1 U18 ( .IN1(n15), .IN2(A[18]), .Q(n16) );
  AND2X1 U19 ( .IN1(n16), .IN2(A[19]), .Q(n17) );
  AND2X1 U20 ( .IN1(n17), .IN2(A[20]), .Q(n18) );
  AND2X1 U21 ( .IN1(n18), .IN2(A[21]), .Q(n19) );
  AND2X1 U22 ( .IN1(n19), .IN2(A[22]), .Q(n20) );
  AND2X1 U23 ( .IN1(n20), .IN2(A[23]), .Q(n21) );
  AND2X1 U24 ( .IN1(n21), .IN2(A[24]), .Q(n22) );
  AND2X1 U25 ( .IN1(n22), .IN2(A[25]), .Q(n23) );
  AND2X1 U26 ( .IN1(n23), .IN2(A[26]), .Q(n24) );
  AND2X1 U27 ( .IN1(n24), .IN2(A[27]), .Q(n25) );
  AND2X1 U28 ( .IN1(n25), .IN2(A[28]), .Q(n26) );
  AND2X1 U29 ( .IN1(n26), .IN2(A[29]), .Q(n27) );
  INVX0 U30 ( .INP(A[2]), .ZN(SUM[2]) );
  XOR2X1 U31 ( .IN1(n27), .IN2(A[30]), .Q(SUM[30]) );
  XOR2X1 U32 ( .IN1(n26), .IN2(A[29]), .Q(SUM[29]) );
  XOR2X1 U33 ( .IN1(n25), .IN2(A[28]), .Q(SUM[28]) );
  XOR2X1 U34 ( .IN1(n24), .IN2(A[27]), .Q(SUM[27]) );
  XOR2X1 U35 ( .IN1(n23), .IN2(A[26]), .Q(SUM[26]) );
  XOR2X1 U36 ( .IN1(n22), .IN2(A[25]), .Q(SUM[25]) );
  XOR2X1 U37 ( .IN1(n21), .IN2(A[24]), .Q(SUM[24]) );
  XOR2X1 U38 ( .IN1(n20), .IN2(A[23]), .Q(SUM[23]) );
  XOR2X1 U39 ( .IN1(n19), .IN2(A[22]), .Q(SUM[22]) );
  XOR2X1 U40 ( .IN1(n18), .IN2(A[21]), .Q(SUM[21]) );
  XOR2X1 U41 ( .IN1(n17), .IN2(A[20]), .Q(SUM[20]) );
  XOR2X1 U42 ( .IN1(n16), .IN2(A[19]), .Q(SUM[19]) );
  XOR2X1 U43 ( .IN1(n15), .IN2(A[18]), .Q(SUM[18]) );
  XOR2X1 U44 ( .IN1(n14), .IN2(A[17]), .Q(SUM[17]) );
  XOR2X1 U45 ( .IN1(n13), .IN2(A[16]), .Q(SUM[16]) );
  XOR2X1 U46 ( .IN1(n12), .IN2(A[15]), .Q(SUM[15]) );
  XOR2X1 U47 ( .IN1(n11), .IN2(A[14]), .Q(SUM[14]) );
  XOR2X1 U48 ( .IN1(n10), .IN2(A[13]), .Q(SUM[13]) );
  XOR2X1 U49 ( .IN1(n9), .IN2(A[12]), .Q(SUM[12]) );
  XOR2X1 U50 ( .IN1(n8), .IN2(A[11]), .Q(SUM[11]) );
  XOR2X1 U51 ( .IN1(n7), .IN2(A[10]), .Q(SUM[10]) );
  XOR2X1 U52 ( .IN1(n6), .IN2(A[9]), .Q(SUM[9]) );
  XOR2X1 U53 ( .IN1(n5), .IN2(A[8]), .Q(SUM[8]) );
  XOR2X1 U54 ( .IN1(n4), .IN2(A[7]), .Q(SUM[7]) );
  XOR2X1 U55 ( .IN1(n3), .IN2(A[6]), .Q(SUM[6]) );
  XOR2X1 U56 ( .IN1(n2), .IN2(A[5]), .Q(SUM[5]) );
  XOR2X1 U57 ( .IN1(n1), .IN2(A[4]), .Q(SUM[4]) );
  XOR2X1 U58 ( .IN1(A[2]), .IN2(A[3]), .Q(SUM[3]) );
endmodule


module pipeline_riscv ( clk, nrst, inst, data_in, inst_addr, data_addr, 
        data_out, data_wr, pc_IF, pc_ID, pc_EXE, pc_MEM, pc_WB );
  input [31:0] inst;
  input [31:0] data_in;
  output [31:0] inst_addr;
  output [31:0] data_addr;
  output [31:0] data_out;
  output [31:0] pc_IF;
  output [31:0] pc_ID;
  output [31:0] pc_EXE;
  output [31:0] pc_MEM;
  output [31:0] pc_WB;
  input clk, nrst;
  output data_wr;
  wire   stall, jal, jr, sw, use_imm, wr_rf, zero, load, jal_pc, n24, n25, n26,
         n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n105, n106, n107, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330;
  wire   [31:0] pc_p4_IF;
  wire   [2:0] sel_pc;
  wire   [31:0] next_pc;
  wire   [31:0] bra_pc;
  wire   [13:9] imm_j;
  wire   [2:0] fwd_jr;
  wire   [31:0] fwd0;
  wire   [4:0] rd;
  wire   [4:0] rs1;
  wire   [4:0] rs2;
  wire   [6:0] funct;
  wire   [8:0] imm_alu;
  wire   [31:0] opA_ID;
  wire   [31:0] opB_ID;
  wire   [31:0] pc_p4_ID;
  wire   [31:0] mem_data_ID;
  wire   [4:0] reg_addr_ID;
  wire   [1:0] flush;
  wire   [4:0] reg_addr_WB;
  wire   [31:0] reg_data_WB;
  wire   [31:0] pc_p4_EXE;
  wire   [31:0] bra_off_EXE;
  wire   [2:0] fwd_opA;
  wire   [31:0] opA;
  wire   [31:0] fwd3;
  wire   [31:0] opA_EXE;
  wire   [2:0] fwd_opB;
  wire   [31:0] opB;
  wire   [31:0] opB_EXE;
  wire   [2:0] fwd_sw;
  wire   [31:0] mem_data_EXE;
  wire   [31:0] mem_data_EXE0;
  wire   [4:0] reg_addr_EXE;
  wire   [6:0] alu_code;
  wire   [31:0] reg_data_MEM;
  wire   [31:0] pc_p4_MEM;
  wire   [4:0] reg_addr_MEM;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133;
  assign inst_addr[31] = pc_IF[31];
  assign inst_addr[30] = pc_IF[30];
  assign inst_addr[29] = pc_IF[29];
  assign inst_addr[28] = pc_IF[28];
  assign inst_addr[27] = pc_IF[27];
  assign inst_addr[26] = pc_IF[26];
  assign inst_addr[25] = pc_IF[25];
  assign inst_addr[24] = pc_IF[24];
  assign inst_addr[23] = pc_IF[23];
  assign inst_addr[22] = pc_IF[22];
  assign inst_addr[21] = pc_IF[21];
  assign inst_addr[20] = pc_IF[20];
  assign inst_addr[19] = pc_IF[19];
  assign inst_addr[18] = pc_IF[18];
  assign inst_addr[17] = pc_IF[17];
  assign inst_addr[16] = pc_IF[16];
  assign inst_addr[15] = pc_IF[15];
  assign inst_addr[14] = pc_IF[14];
  assign inst_addr[13] = pc_IF[13];
  assign inst_addr[12] = pc_IF[12];
  assign inst_addr[11] = pc_IF[11];
  assign inst_addr[10] = pc_IF[10];
  assign inst_addr[9] = pc_IF[9];
  assign inst_addr[8] = pc_IF[8];
  assign inst_addr[7] = pc_IF[7];
  assign inst_addr[6] = pc_IF[6];
  assign inst_addr[5] = pc_IF[5];
  assign inst_addr[4] = pc_IF[4];
  assign inst_addr[3] = pc_IF[3];
  assign inst_addr[2] = pc_IF[2];
  assign inst_addr[1] = pc_IF[1];
  assign inst_addr[0] = pc_IF[0];

  AO22X1 U91 ( .IN1(rd[4]), .IN2(n322), .IN3(imm_alu[8]), .IN4(n24), .Q(rs2[4]) );
  AO22X1 U92 ( .IN1(rd[3]), .IN2(n322), .IN3(imm_alu[7]), .IN4(n24), .Q(rs2[3]) );
  AO22X1 U93 ( .IN1(rd[2]), .IN2(n322), .IN3(imm_alu[6]), .IN4(n24), .Q(rs2[2]) );
  AO22X1 U94 ( .IN1(rd[1]), .IN2(n322), .IN3(imm_alu[5]), .IN4(n24), .Q(rs2[1]) );
  AO22X1 U95 ( .IN1(rd[0]), .IN2(n322), .IN3(imm_alu[4]), .IN4(n24), .Q(rs2[0]) );
  AND2X1 U96 ( .IN1(n316), .IN2(imm_j[13]), .Q(rs1[4]) );
  AND2X1 U97 ( .IN1(n316), .IN2(imm_j[12]), .Q(rs1[3]) );
  AND2X1 U98 ( .IN1(n316), .IN2(imm_j[11]), .Q(rs1[2]) );
  AND2X1 U99 ( .IN1(n316), .IN2(imm_j[10]), .Q(rs1[1]) );
  AND2X1 U100 ( .IN1(n316), .IN2(imm_j[9]), .Q(rs1[0]) );
  AO222X1 U101 ( .IN1(pc_p4_MEM[9]), .IN2(n25), .IN3(data_addr[9]), .IN4(n286), 
        .IN5(load), .IN6(data_in[9]), .Q(reg_data_MEM[9]) );
  AO222X1 U102 ( .IN1(pc_p4_MEM[8]), .IN2(n284), .IN3(data_addr[8]), .IN4(n285), .IN5(data_in[8]), .IN6(load), .Q(reg_data_MEM[8]) );
  AO222X1 U103 ( .IN1(pc_p4_MEM[7]), .IN2(n25), .IN3(data_addr[7]), .IN4(n26), 
        .IN5(data_in[7]), .IN6(load), .Q(reg_data_MEM[7]) );
  AO222X1 U104 ( .IN1(pc_p4_MEM[6]), .IN2(n284), .IN3(data_addr[6]), .IN4(n286), .IN5(data_in[6]), .IN6(load), .Q(reg_data_MEM[6]) );
  AO222X1 U105 ( .IN1(pc_p4_MEM[5]), .IN2(n25), .IN3(data_addr[5]), .IN4(n285), 
        .IN5(data_in[5]), .IN6(load), .Q(reg_data_MEM[5]) );
  AO222X1 U106 ( .IN1(pc_p4_MEM[4]), .IN2(n284), .IN3(data_addr[4]), .IN4(n26), 
        .IN5(data_in[4]), .IN6(load), .Q(reg_data_MEM[4]) );
  AO222X1 U107 ( .IN1(pc_p4_MEM[3]), .IN2(n25), .IN3(data_addr[3]), .IN4(n286), 
        .IN5(data_in[3]), .IN6(load), .Q(reg_data_MEM[3]) );
  AO222X1 U108 ( .IN1(pc_p4_MEM[31]), .IN2(n284), .IN3(data_addr[31]), .IN4(
        n285), .IN5(data_in[31]), .IN6(load), .Q(reg_data_MEM[31]) );
  AO222X1 U109 ( .IN1(pc_p4_MEM[30]), .IN2(n25), .IN3(data_addr[30]), .IN4(n26), .IN5(data_in[30]), .IN6(load), .Q(reg_data_MEM[30]) );
  AO222X1 U110 ( .IN1(pc_p4_MEM[2]), .IN2(n284), .IN3(data_addr[2]), .IN4(n286), .IN5(data_in[2]), .IN6(load), .Q(reg_data_MEM[2]) );
  AO222X1 U111 ( .IN1(pc_p4_MEM[29]), .IN2(n25), .IN3(data_addr[29]), .IN4(
        n285), .IN5(data_in[29]), .IN6(load), .Q(reg_data_MEM[29]) );
  AO222X1 U112 ( .IN1(pc_p4_MEM[28]), .IN2(n284), .IN3(data_addr[28]), .IN4(
        n26), .IN5(data_in[28]), .IN6(load), .Q(reg_data_MEM[28]) );
  AO222X1 U113 ( .IN1(pc_p4_MEM[27]), .IN2(n25), .IN3(data_addr[27]), .IN4(
        n286), .IN5(data_in[27]), .IN6(load), .Q(reg_data_MEM[27]) );
  AO222X1 U114 ( .IN1(pc_p4_MEM[26]), .IN2(n284), .IN3(data_addr[26]), .IN4(
        n285), .IN5(data_in[26]), .IN6(load), .Q(reg_data_MEM[26]) );
  AO222X1 U115 ( .IN1(pc_p4_MEM[25]), .IN2(n25), .IN3(data_addr[25]), .IN4(n26), .IN5(data_in[25]), .IN6(load), .Q(reg_data_MEM[25]) );
  AO222X1 U116 ( .IN1(pc_p4_MEM[24]), .IN2(n284), .IN3(data_addr[24]), .IN4(
        n286), .IN5(data_in[24]), .IN6(load), .Q(reg_data_MEM[24]) );
  AO222X1 U117 ( .IN1(pc_p4_MEM[23]), .IN2(n25), .IN3(data_addr[23]), .IN4(
        n285), .IN5(data_in[23]), .IN6(load), .Q(reg_data_MEM[23]) );
  AO222X1 U118 ( .IN1(pc_p4_MEM[22]), .IN2(n284), .IN3(data_addr[22]), .IN4(
        n26), .IN5(data_in[22]), .IN6(load), .Q(reg_data_MEM[22]) );
  AO222X1 U119 ( .IN1(pc_p4_MEM[21]), .IN2(n25), .IN3(data_addr[21]), .IN4(
        n286), .IN5(data_in[21]), .IN6(load), .Q(reg_data_MEM[21]) );
  AO222X1 U120 ( .IN1(pc_p4_MEM[20]), .IN2(n284), .IN3(data_addr[20]), .IN4(
        n285), .IN5(data_in[20]), .IN6(load), .Q(reg_data_MEM[20]) );
  AO222X1 U121 ( .IN1(pc_p4_MEM[1]), .IN2(n25), .IN3(data_addr[1]), .IN4(n26), 
        .IN5(data_in[1]), .IN6(load), .Q(reg_data_MEM[1]) );
  AO222X1 U122 ( .IN1(pc_p4_MEM[19]), .IN2(n284), .IN3(data_addr[19]), .IN4(
        n286), .IN5(data_in[19]), .IN6(load), .Q(reg_data_MEM[19]) );
  AO222X1 U123 ( .IN1(pc_p4_MEM[18]), .IN2(n25), .IN3(data_addr[18]), .IN4(
        n285), .IN5(data_in[18]), .IN6(load), .Q(reg_data_MEM[18]) );
  AO222X1 U124 ( .IN1(pc_p4_MEM[17]), .IN2(n284), .IN3(data_addr[17]), .IN4(
        n26), .IN5(data_in[17]), .IN6(load), .Q(reg_data_MEM[17]) );
  AO222X1 U125 ( .IN1(pc_p4_MEM[16]), .IN2(n25), .IN3(data_addr[16]), .IN4(
        n286), .IN5(data_in[16]), .IN6(load), .Q(reg_data_MEM[16]) );
  AO222X1 U126 ( .IN1(pc_p4_MEM[15]), .IN2(n284), .IN3(data_addr[15]), .IN4(
        n285), .IN5(data_in[15]), .IN6(load), .Q(reg_data_MEM[15]) );
  AO222X1 U127 ( .IN1(pc_p4_MEM[14]), .IN2(n25), .IN3(data_addr[14]), .IN4(n26), .IN5(data_in[14]), .IN6(load), .Q(reg_data_MEM[14]) );
  AO222X1 U128 ( .IN1(pc_p4_MEM[13]), .IN2(n284), .IN3(data_addr[13]), .IN4(
        n286), .IN5(data_in[13]), .IN6(load), .Q(reg_data_MEM[13]) );
  AO222X1 U129 ( .IN1(pc_p4_MEM[12]), .IN2(n25), .IN3(data_addr[12]), .IN4(
        n285), .IN5(data_in[12]), .IN6(load), .Q(reg_data_MEM[12]) );
  AO222X1 U130 ( .IN1(pc_p4_MEM[11]), .IN2(n284), .IN3(data_addr[11]), .IN4(
        n26), .IN5(data_in[11]), .IN6(load), .Q(reg_data_MEM[11]) );
  AO222X1 U131 ( .IN1(pc_p4_MEM[10]), .IN2(n25), .IN3(data_addr[10]), .IN4(
        n286), .IN5(data_in[10]), .IN6(load), .Q(reg_data_MEM[10]) );
  AO222X1 U132 ( .IN1(pc_p4_MEM[0]), .IN2(n284), .IN3(data_addr[0]), .IN4(n285), .IN5(data_in[0]), .IN6(load), .Q(reg_data_MEM[0]) );
  AND2X1 U133 ( .IN1(n316), .IN2(rd[4]), .Q(reg_addr_ID[4]) );
  AND2X1 U134 ( .IN1(n316), .IN2(rd[3]), .Q(reg_addr_ID[3]) );
  AND2X1 U135 ( .IN1(n316), .IN2(rd[2]), .Q(reg_addr_ID[2]) );
  AND2X1 U136 ( .IN1(n316), .IN2(rd[1]), .Q(reg_addr_ID[1]) );
  OR2X1 U137 ( .IN1(rd[0]), .IN2(n314), .Q(reg_addr_ID[0]) );
  AO222X1 U138 ( .IN1(funct[0]), .IN2(n27), .IN3(mem_data_ID[9]), .IN4(n28), 
        .IN5(pc_p4_ID[9]), .IN6(n314), .Q(opB_ID[9]) );
  AO222X1 U139 ( .IN1(n27), .IN2(imm_alu[8]), .IN3(mem_data_ID[8]), .IN4(n283), 
        .IN5(pc_p4_ID[8]), .IN6(n315), .Q(opB_ID[8]) );
  AO222X1 U140 ( .IN1(n27), .IN2(imm_alu[7]), .IN3(mem_data_ID[7]), .IN4(n28), 
        .IN5(pc_p4_ID[7]), .IN6(n315), .Q(opB_ID[7]) );
  AO222X1 U141 ( .IN1(n27), .IN2(imm_alu[6]), .IN3(mem_data_ID[6]), .IN4(n283), 
        .IN5(pc_p4_ID[6]), .IN6(n315), .Q(opB_ID[6]) );
  AO222X1 U142 ( .IN1(n27), .IN2(imm_alu[5]), .IN3(mem_data_ID[5]), .IN4(n28), 
        .IN5(pc_p4_ID[5]), .IN6(n315), .Q(opB_ID[5]) );
  AO222X1 U143 ( .IN1(n27), .IN2(imm_alu[4]), .IN3(mem_data_ID[4]), .IN4(n283), 
        .IN5(pc_p4_ID[4]), .IN6(n314), .Q(opB_ID[4]) );
  AO222X1 U144 ( .IN1(imm_alu[3]), .IN2(n27), .IN3(mem_data_ID[3]), .IN4(n28), 
        .IN5(pc_p4_ID[3]), .IN6(n314), .Q(opB_ID[3]) );
  AO221X1 U145 ( .IN1(mem_data_ID[31]), .IN2(n283), .IN3(pc_p4_ID[31]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[31]) );
  AO221X1 U146 ( .IN1(mem_data_ID[30]), .IN2(n28), .IN3(pc_p4_ID[30]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[30]) );
  AO222X1 U147 ( .IN1(imm_alu[2]), .IN2(n27), .IN3(mem_data_ID[2]), .IN4(n283), 
        .IN5(pc_p4_ID[2]), .IN6(n314), .Q(opB_ID[2]) );
  AO221X1 U148 ( .IN1(mem_data_ID[29]), .IN2(n283), .IN3(pc_p4_ID[29]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[29]) );
  AO221X1 U149 ( .IN1(mem_data_ID[28]), .IN2(n28), .IN3(pc_p4_ID[28]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[28]) );
  AO221X1 U150 ( .IN1(mem_data_ID[27]), .IN2(n283), .IN3(pc_p4_ID[27]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[27]) );
  AO221X1 U151 ( .IN1(mem_data_ID[26]), .IN2(n28), .IN3(pc_p4_ID[26]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[26]) );
  AO221X1 U152 ( .IN1(mem_data_ID[25]), .IN2(n283), .IN3(pc_p4_ID[25]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[25]) );
  AO221X1 U153 ( .IN1(mem_data_ID[24]), .IN2(n28), .IN3(pc_p4_ID[24]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[24]) );
  AO221X1 U154 ( .IN1(mem_data_ID[23]), .IN2(n283), .IN3(pc_p4_ID[23]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[23]) );
  AO221X1 U155 ( .IN1(mem_data_ID[22]), .IN2(n28), .IN3(pc_p4_ID[22]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[22]) );
  AO221X1 U156 ( .IN1(mem_data_ID[21]), .IN2(n283), .IN3(pc_p4_ID[21]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[21]) );
  AO221X1 U157 ( .IN1(mem_data_ID[20]), .IN2(n28), .IN3(pc_p4_ID[20]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[20]) );
  AO222X1 U158 ( .IN1(imm_alu[1]), .IN2(n27), .IN3(mem_data_ID[1]), .IN4(n28), 
        .IN5(pc_p4_ID[1]), .IN6(n314), .Q(opB_ID[1]) );
  AO221X1 U159 ( .IN1(mem_data_ID[19]), .IN2(n283), .IN3(pc_p4_ID[19]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[19]) );
  AO221X1 U160 ( .IN1(mem_data_ID[18]), .IN2(n28), .IN3(pc_p4_ID[18]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[18]) );
  AO221X1 U161 ( .IN1(mem_data_ID[17]), .IN2(n283), .IN3(pc_p4_ID[17]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[17]) );
  AO221X1 U162 ( .IN1(mem_data_ID[16]), .IN2(n28), .IN3(pc_p4_ID[16]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[16]) );
  AO221X1 U163 ( .IN1(mem_data_ID[15]), .IN2(n283), .IN3(pc_p4_ID[15]), .IN4(
        n314), .IN5(n29), .Q(opB_ID[15]) );
  AO222X1 U165 ( .IN1(funct[5]), .IN2(n27), .IN3(mem_data_ID[14]), .IN4(n283), 
        .IN5(pc_p4_ID[14]), .IN6(n314), .Q(opB_ID[14]) );
  AO222X1 U166 ( .IN1(funct[4]), .IN2(n27), .IN3(mem_data_ID[13]), .IN4(n28), 
        .IN5(pc_p4_ID[13]), .IN6(n314), .Q(opB_ID[13]) );
  AO222X1 U167 ( .IN1(funct[3]), .IN2(n27), .IN3(mem_data_ID[12]), .IN4(n283), 
        .IN5(pc_p4_ID[12]), .IN6(n314), .Q(opB_ID[12]) );
  AO222X1 U168 ( .IN1(funct[2]), .IN2(n27), .IN3(mem_data_ID[11]), .IN4(n28), 
        .IN5(pc_p4_ID[11]), .IN6(n314), .Q(opB_ID[11]) );
  AO222X1 U169 ( .IN1(funct[1]), .IN2(n27), .IN3(mem_data_ID[10]), .IN4(n283), 
        .IN5(pc_p4_ID[10]), .IN6(n314), .Q(opB_ID[10]) );
  AO222X1 U170 ( .IN1(imm_alu[0]), .IN2(n27), .IN3(mem_data_ID[0]), .IN4(n28), 
        .IN5(pc_p4_ID[0]), .IN6(n314), .Q(opB_ID[0]) );
  AO221X1 U172 ( .IN1(opB_EXE[9]), .IN2(n311), .IN3(fwd3[9]), .IN4(n308), 
        .IN5(n32), .Q(opB[9]) );
  AO22X1 U173 ( .IN1(fwd_opB[2]), .IN2(data_addr[9]), .IN3(reg_data_WB[9]), 
        .IN4(n282), .Q(n32) );
  AO221X1 U174 ( .IN1(opB_EXE[8]), .IN2(n311), .IN3(fwd3[8]), .IN4(n308), 
        .IN5(n34), .Q(opB[8]) );
  AO22X1 U175 ( .IN1(fwd_opB[2]), .IN2(data_addr[8]), .IN3(reg_data_WB[8]), 
        .IN4(n281), .Q(n34) );
  AO221X1 U176 ( .IN1(opB_EXE[7]), .IN2(n311), .IN3(fwd3[7]), .IN4(n308), 
        .IN5(n35), .Q(opB[7]) );
  AO22X1 U177 ( .IN1(fwd_opB[2]), .IN2(data_addr[7]), .IN3(reg_data_WB[7]), 
        .IN4(n33), .Q(n35) );
  AO221X1 U178 ( .IN1(opB_EXE[6]), .IN2(n311), .IN3(fwd3[6]), .IN4(n308), 
        .IN5(n36), .Q(opB[6]) );
  AO22X1 U179 ( .IN1(fwd_opB[2]), .IN2(data_addr[6]), .IN3(reg_data_WB[6]), 
        .IN4(n282), .Q(n36) );
  AO221X1 U180 ( .IN1(opB_EXE[5]), .IN2(n311), .IN3(fwd3[5]), .IN4(n308), 
        .IN5(n37), .Q(opB[5]) );
  AO22X1 U181 ( .IN1(fwd_opB[2]), .IN2(data_addr[5]), .IN3(reg_data_WB[5]), 
        .IN4(n281), .Q(n37) );
  AO221X1 U182 ( .IN1(opB_EXE[4]), .IN2(n311), .IN3(fwd3[4]), .IN4(n308), 
        .IN5(n38), .Q(opB[4]) );
  AO22X1 U183 ( .IN1(fwd_opB[2]), .IN2(data_addr[4]), .IN3(reg_data_WB[4]), 
        .IN4(n33), .Q(n38) );
  AO221X1 U184 ( .IN1(opB_EXE[3]), .IN2(n311), .IN3(fwd3[3]), .IN4(n308), 
        .IN5(n39), .Q(opB[3]) );
  AO22X1 U185 ( .IN1(fwd_opB[2]), .IN2(data_addr[3]), .IN3(reg_data_WB[3]), 
        .IN4(n282), .Q(n39) );
  AO221X1 U186 ( .IN1(opB_EXE[31]), .IN2(n311), .IN3(fwd3[31]), .IN4(n308), 
        .IN5(n40), .Q(opB[31]) );
  AO22X1 U187 ( .IN1(fwd_opB[2]), .IN2(data_addr[31]), .IN3(reg_data_WB[31]), 
        .IN4(n281), .Q(n40) );
  AO221X1 U188 ( .IN1(opB_EXE[30]), .IN2(n311), .IN3(fwd3[30]), .IN4(n308), 
        .IN5(n41), .Q(opB[30]) );
  AO22X1 U189 ( .IN1(fwd_opB[2]), .IN2(data_addr[30]), .IN3(reg_data_WB[30]), 
        .IN4(n33), .Q(n41) );
  AO221X1 U190 ( .IN1(opB_EXE[2]), .IN2(n311), .IN3(fwd3[2]), .IN4(n308), 
        .IN5(n42), .Q(opB[2]) );
  AO22X1 U191 ( .IN1(fwd_opB[2]), .IN2(data_addr[2]), .IN3(reg_data_WB[2]), 
        .IN4(n282), .Q(n42) );
  AO221X1 U192 ( .IN1(opB_EXE[29]), .IN2(n311), .IN3(fwd3[29]), .IN4(n308), 
        .IN5(n43), .Q(opB[29]) );
  AO22X1 U193 ( .IN1(fwd_opB[2]), .IN2(data_addr[29]), .IN3(reg_data_WB[29]), 
        .IN4(n281), .Q(n43) );
  AO221X1 U194 ( .IN1(opB_EXE[28]), .IN2(n311), .IN3(fwd3[28]), .IN4(n308), 
        .IN5(n44), .Q(opB[28]) );
  AO22X1 U195 ( .IN1(fwd_opB[2]), .IN2(data_addr[28]), .IN3(reg_data_WB[28]), 
        .IN4(n33), .Q(n44) );
  AO221X1 U196 ( .IN1(opB_EXE[27]), .IN2(n312), .IN3(fwd3[27]), .IN4(n309), 
        .IN5(n45), .Q(opB[27]) );
  AO22X1 U197 ( .IN1(fwd_opB[2]), .IN2(data_addr[27]), .IN3(reg_data_WB[27]), 
        .IN4(n282), .Q(n45) );
  AO221X1 U198 ( .IN1(opB_EXE[26]), .IN2(n312), .IN3(fwd3[26]), .IN4(n309), 
        .IN5(n46), .Q(opB[26]) );
  AO22X1 U199 ( .IN1(fwd_opB[2]), .IN2(data_addr[26]), .IN3(reg_data_WB[26]), 
        .IN4(n281), .Q(n46) );
  AO221X1 U200 ( .IN1(opB_EXE[25]), .IN2(n312), .IN3(fwd3[25]), .IN4(n309), 
        .IN5(n47), .Q(opB[25]) );
  AO22X1 U201 ( .IN1(fwd_opB[2]), .IN2(data_addr[25]), .IN3(reg_data_WB[25]), 
        .IN4(n33), .Q(n47) );
  AO221X1 U202 ( .IN1(opB_EXE[24]), .IN2(n312), .IN3(fwd3[24]), .IN4(n309), 
        .IN5(n48), .Q(opB[24]) );
  AO22X1 U203 ( .IN1(fwd_opB[2]), .IN2(data_addr[24]), .IN3(reg_data_WB[24]), 
        .IN4(n282), .Q(n48) );
  AO221X1 U204 ( .IN1(opB_EXE[23]), .IN2(n312), .IN3(fwd3[23]), .IN4(n309), 
        .IN5(n49), .Q(opB[23]) );
  AO22X1 U205 ( .IN1(fwd_opB[2]), .IN2(data_addr[23]), .IN3(reg_data_WB[23]), 
        .IN4(n281), .Q(n49) );
  AO221X1 U206 ( .IN1(opB_EXE[22]), .IN2(n312), .IN3(fwd3[22]), .IN4(n309), 
        .IN5(n50), .Q(opB[22]) );
  AO22X1 U207 ( .IN1(fwd_opB[2]), .IN2(data_addr[22]), .IN3(reg_data_WB[22]), 
        .IN4(n33), .Q(n50) );
  AO221X1 U208 ( .IN1(opB_EXE[21]), .IN2(n312), .IN3(fwd3[21]), .IN4(n309), 
        .IN5(n51), .Q(opB[21]) );
  AO22X1 U209 ( .IN1(fwd_opB[2]), .IN2(data_addr[21]), .IN3(reg_data_WB[21]), 
        .IN4(n282), .Q(n51) );
  AO221X1 U210 ( .IN1(opB_EXE[20]), .IN2(n312), .IN3(fwd3[20]), .IN4(n309), 
        .IN5(n52), .Q(opB[20]) );
  AO22X1 U211 ( .IN1(fwd_opB[2]), .IN2(data_addr[20]), .IN3(reg_data_WB[20]), 
        .IN4(n281), .Q(n52) );
  AO221X1 U212 ( .IN1(opB_EXE[1]), .IN2(n312), .IN3(fwd3[1]), .IN4(n309), 
        .IN5(n53), .Q(opB[1]) );
  AO22X1 U213 ( .IN1(fwd_opB[2]), .IN2(data_addr[1]), .IN3(reg_data_WB[1]), 
        .IN4(n33), .Q(n53) );
  AO221X1 U214 ( .IN1(opB_EXE[19]), .IN2(n312), .IN3(fwd3[19]), .IN4(n309), 
        .IN5(n54), .Q(opB[19]) );
  AO22X1 U215 ( .IN1(fwd_opB[2]), .IN2(data_addr[19]), .IN3(reg_data_WB[19]), 
        .IN4(n282), .Q(n54) );
  AO221X1 U216 ( .IN1(opB_EXE[18]), .IN2(n312), .IN3(fwd3[18]), .IN4(n309), 
        .IN5(n55), .Q(opB[18]) );
  AO22X1 U217 ( .IN1(fwd_opB[2]), .IN2(data_addr[18]), .IN3(reg_data_WB[18]), 
        .IN4(n281), .Q(n55) );
  AO221X1 U218 ( .IN1(opB_EXE[17]), .IN2(n312), .IN3(fwd3[17]), .IN4(n309), 
        .IN5(n56), .Q(opB[17]) );
  AO22X1 U219 ( .IN1(fwd_opB[2]), .IN2(data_addr[17]), .IN3(reg_data_WB[17]), 
        .IN4(n33), .Q(n56) );
  AO221X1 U220 ( .IN1(opB_EXE[16]), .IN2(n313), .IN3(fwd3[16]), .IN4(n310), 
        .IN5(n57), .Q(opB[16]) );
  AO22X1 U221 ( .IN1(fwd_opB[2]), .IN2(data_addr[16]), .IN3(reg_data_WB[16]), 
        .IN4(n282), .Q(n57) );
  AO221X1 U222 ( .IN1(opB_EXE[15]), .IN2(n313), .IN3(fwd3[15]), .IN4(n310), 
        .IN5(n58), .Q(opB[15]) );
  AO22X1 U223 ( .IN1(fwd_opB[2]), .IN2(data_addr[15]), .IN3(reg_data_WB[15]), 
        .IN4(n281), .Q(n58) );
  AO221X1 U224 ( .IN1(opB_EXE[14]), .IN2(n313), .IN3(fwd3[14]), .IN4(n310), 
        .IN5(n59), .Q(opB[14]) );
  AO22X1 U225 ( .IN1(fwd_opB[2]), .IN2(data_addr[14]), .IN3(reg_data_WB[14]), 
        .IN4(n33), .Q(n59) );
  AO221X1 U226 ( .IN1(opB_EXE[13]), .IN2(n313), .IN3(fwd3[13]), .IN4(n310), 
        .IN5(n60), .Q(opB[13]) );
  AO22X1 U227 ( .IN1(fwd_opB[2]), .IN2(data_addr[13]), .IN3(reg_data_WB[13]), 
        .IN4(n282), .Q(n60) );
  AO221X1 U228 ( .IN1(opB_EXE[12]), .IN2(n313), .IN3(fwd3[12]), .IN4(n310), 
        .IN5(n61), .Q(opB[12]) );
  AO22X1 U229 ( .IN1(fwd_opB[2]), .IN2(data_addr[12]), .IN3(reg_data_WB[12]), 
        .IN4(n281), .Q(n61) );
  AO221X1 U230 ( .IN1(opB_EXE[11]), .IN2(n313), .IN3(fwd3[11]), .IN4(n310), 
        .IN5(n62), .Q(opB[11]) );
  AO22X1 U231 ( .IN1(fwd_opB[2]), .IN2(data_addr[11]), .IN3(reg_data_WB[11]), 
        .IN4(n33), .Q(n62) );
  AO221X1 U232 ( .IN1(opB_EXE[10]), .IN2(n313), .IN3(fwd3[10]), .IN4(n310), 
        .IN5(n63), .Q(opB[10]) );
  AO22X1 U233 ( .IN1(fwd_opB[2]), .IN2(data_addr[10]), .IN3(reg_data_WB[10]), 
        .IN4(n282), .Q(n63) );
  AO221X1 U234 ( .IN1(opB_EXE[0]), .IN2(n313), .IN3(fwd3[0]), .IN4(n310), 
        .IN5(n64), .Q(opB[0]) );
  AO22X1 U235 ( .IN1(fwd_opB[2]), .IN2(data_addr[0]), .IN3(reg_data_WB[0]), 
        .IN4(n281), .Q(n64) );
  AO221X1 U238 ( .IN1(opA_EXE[9]), .IN2(n305), .IN3(n302), .IN4(fwd3[9]), 
        .IN5(n67), .Q(opA[9]) );
  AO22X1 U239 ( .IN1(fwd_opA[2]), .IN2(data_addr[9]), .IN3(n280), .IN4(
        reg_data_WB[9]), .Q(n67) );
  AO221X1 U240 ( .IN1(opA_EXE[8]), .IN2(n305), .IN3(n302), .IN4(fwd3[8]), 
        .IN5(n69), .Q(opA[8]) );
  AO22X1 U241 ( .IN1(fwd_opA[2]), .IN2(data_addr[8]), .IN3(n279), .IN4(
        reg_data_WB[8]), .Q(n69) );
  AO221X1 U242 ( .IN1(opA_EXE[7]), .IN2(n305), .IN3(n302), .IN4(fwd3[7]), 
        .IN5(n70), .Q(opA[7]) );
  AO22X1 U243 ( .IN1(fwd_opA[2]), .IN2(data_addr[7]), .IN3(n68), .IN4(
        reg_data_WB[7]), .Q(n70) );
  AO221X1 U244 ( .IN1(opA_EXE[6]), .IN2(n305), .IN3(n302), .IN4(fwd3[6]), 
        .IN5(n71), .Q(opA[6]) );
  AO22X1 U245 ( .IN1(fwd_opA[2]), .IN2(data_addr[6]), .IN3(n280), .IN4(
        reg_data_WB[6]), .Q(n71) );
  AO221X1 U246 ( .IN1(opA_EXE[5]), .IN2(n305), .IN3(n302), .IN4(fwd3[5]), 
        .IN5(n72), .Q(opA[5]) );
  AO22X1 U247 ( .IN1(fwd_opA[2]), .IN2(data_addr[5]), .IN3(n279), .IN4(
        reg_data_WB[5]), .Q(n72) );
  AO221X1 U248 ( .IN1(opA_EXE[4]), .IN2(n305), .IN3(n302), .IN4(fwd3[4]), 
        .IN5(n73), .Q(opA[4]) );
  AO22X1 U249 ( .IN1(fwd_opA[2]), .IN2(data_addr[4]), .IN3(n68), .IN4(
        reg_data_WB[4]), .Q(n73) );
  AO221X1 U250 ( .IN1(opA_EXE[3]), .IN2(n305), .IN3(n302), .IN4(fwd3[3]), 
        .IN5(n74), .Q(opA[3]) );
  AO22X1 U251 ( .IN1(fwd_opA[2]), .IN2(data_addr[3]), .IN3(n280), .IN4(
        reg_data_WB[3]), .Q(n74) );
  AO221X1 U252 ( .IN1(opA_EXE[31]), .IN2(n305), .IN3(n302), .IN4(fwd3[31]), 
        .IN5(n75), .Q(opA[31]) );
  AO22X1 U253 ( .IN1(fwd_opA[2]), .IN2(data_addr[31]), .IN3(n279), .IN4(
        reg_data_WB[31]), .Q(n75) );
  AO221X1 U254 ( .IN1(opA_EXE[30]), .IN2(n305), .IN3(n302), .IN4(fwd3[30]), 
        .IN5(n76), .Q(opA[30]) );
  AO22X1 U255 ( .IN1(fwd_opA[2]), .IN2(data_addr[30]), .IN3(n68), .IN4(
        reg_data_WB[30]), .Q(n76) );
  AO221X1 U256 ( .IN1(opA_EXE[2]), .IN2(n305), .IN3(n302), .IN4(fwd3[2]), 
        .IN5(n77), .Q(opA[2]) );
  AO22X1 U257 ( .IN1(fwd_opA[2]), .IN2(data_addr[2]), .IN3(n280), .IN4(
        reg_data_WB[2]), .Q(n77) );
  AO221X1 U258 ( .IN1(opA_EXE[29]), .IN2(n305), .IN3(n302), .IN4(fwd3[29]), 
        .IN5(n78), .Q(opA[29]) );
  AO22X1 U259 ( .IN1(fwd_opA[2]), .IN2(data_addr[29]), .IN3(n279), .IN4(
        reg_data_WB[29]), .Q(n78) );
  AO221X1 U260 ( .IN1(opA_EXE[28]), .IN2(n305), .IN3(n302), .IN4(fwd3[28]), 
        .IN5(n79), .Q(opA[28]) );
  AO22X1 U261 ( .IN1(fwd_opA[2]), .IN2(data_addr[28]), .IN3(n68), .IN4(
        reg_data_WB[28]), .Q(n79) );
  AO221X1 U262 ( .IN1(opA_EXE[27]), .IN2(n306), .IN3(n303), .IN4(fwd3[27]), 
        .IN5(n80), .Q(opA[27]) );
  AO22X1 U263 ( .IN1(fwd_opA[2]), .IN2(data_addr[27]), .IN3(n280), .IN4(
        reg_data_WB[27]), .Q(n80) );
  AO221X1 U264 ( .IN1(opA_EXE[26]), .IN2(n306), .IN3(n303), .IN4(fwd3[26]), 
        .IN5(n81), .Q(opA[26]) );
  AO22X1 U265 ( .IN1(fwd_opA[2]), .IN2(data_addr[26]), .IN3(n279), .IN4(
        reg_data_WB[26]), .Q(n81) );
  AO221X1 U266 ( .IN1(opA_EXE[25]), .IN2(n306), .IN3(n303), .IN4(fwd3[25]), 
        .IN5(n82), .Q(opA[25]) );
  AO22X1 U267 ( .IN1(fwd_opA[2]), .IN2(data_addr[25]), .IN3(n68), .IN4(
        reg_data_WB[25]), .Q(n82) );
  AO221X1 U268 ( .IN1(opA_EXE[24]), .IN2(n306), .IN3(n303), .IN4(fwd3[24]), 
        .IN5(n83), .Q(opA[24]) );
  AO22X1 U269 ( .IN1(fwd_opA[2]), .IN2(data_addr[24]), .IN3(n280), .IN4(
        reg_data_WB[24]), .Q(n83) );
  AO221X1 U270 ( .IN1(opA_EXE[23]), .IN2(n306), .IN3(n303), .IN4(fwd3[23]), 
        .IN5(n84), .Q(opA[23]) );
  AO22X1 U271 ( .IN1(fwd_opA[2]), .IN2(data_addr[23]), .IN3(n279), .IN4(
        reg_data_WB[23]), .Q(n84) );
  AO221X1 U272 ( .IN1(opA_EXE[22]), .IN2(n306), .IN3(n303), .IN4(fwd3[22]), 
        .IN5(n85), .Q(opA[22]) );
  AO22X1 U273 ( .IN1(fwd_opA[2]), .IN2(data_addr[22]), .IN3(n68), .IN4(
        reg_data_WB[22]), .Q(n85) );
  AO221X1 U274 ( .IN1(opA_EXE[21]), .IN2(n306), .IN3(n303), .IN4(fwd3[21]), 
        .IN5(n86), .Q(opA[21]) );
  AO22X1 U275 ( .IN1(fwd_opA[2]), .IN2(data_addr[21]), .IN3(n280), .IN4(
        reg_data_WB[21]), .Q(n86) );
  AO221X1 U276 ( .IN1(opA_EXE[20]), .IN2(n306), .IN3(n303), .IN4(fwd3[20]), 
        .IN5(n87), .Q(opA[20]) );
  AO22X1 U277 ( .IN1(fwd_opA[2]), .IN2(data_addr[20]), .IN3(n279), .IN4(
        reg_data_WB[20]), .Q(n87) );
  AO221X1 U278 ( .IN1(opA_EXE[1]), .IN2(n306), .IN3(n303), .IN4(fwd3[1]), 
        .IN5(n88), .Q(opA[1]) );
  AO22X1 U279 ( .IN1(fwd_opA[2]), .IN2(data_addr[1]), .IN3(n68), .IN4(
        reg_data_WB[1]), .Q(n88) );
  AO221X1 U280 ( .IN1(opA_EXE[19]), .IN2(n306), .IN3(n303), .IN4(fwd3[19]), 
        .IN5(n89), .Q(opA[19]) );
  AO22X1 U281 ( .IN1(fwd_opA[2]), .IN2(data_addr[19]), .IN3(n280), .IN4(
        reg_data_WB[19]), .Q(n89) );
  AO221X1 U282 ( .IN1(opA_EXE[18]), .IN2(n306), .IN3(n303), .IN4(fwd3[18]), 
        .IN5(n90), .Q(opA[18]) );
  AO22X1 U283 ( .IN1(fwd_opA[2]), .IN2(data_addr[18]), .IN3(n279), .IN4(
        reg_data_WB[18]), .Q(n90) );
  AO221X1 U284 ( .IN1(opA_EXE[17]), .IN2(n306), .IN3(n303), .IN4(fwd3[17]), 
        .IN5(n91), .Q(opA[17]) );
  AO22X1 U285 ( .IN1(fwd_opA[2]), .IN2(data_addr[17]), .IN3(n68), .IN4(
        reg_data_WB[17]), .Q(n91) );
  AO221X1 U286 ( .IN1(opA_EXE[16]), .IN2(n307), .IN3(n304), .IN4(fwd3[16]), 
        .IN5(n92), .Q(opA[16]) );
  AO22X1 U287 ( .IN1(fwd_opA[2]), .IN2(data_addr[16]), .IN3(n280), .IN4(
        reg_data_WB[16]), .Q(n92) );
  AO221X1 U288 ( .IN1(opA_EXE[15]), .IN2(n307), .IN3(n304), .IN4(fwd3[15]), 
        .IN5(n93), .Q(opA[15]) );
  AO22X1 U289 ( .IN1(fwd_opA[2]), .IN2(data_addr[15]), .IN3(n279), .IN4(
        reg_data_WB[15]), .Q(n93) );
  AO221X1 U290 ( .IN1(opA_EXE[14]), .IN2(n307), .IN3(n304), .IN4(fwd3[14]), 
        .IN5(n94), .Q(opA[14]) );
  AO22X1 U291 ( .IN1(fwd_opA[2]), .IN2(data_addr[14]), .IN3(n68), .IN4(
        reg_data_WB[14]), .Q(n94) );
  AO221X1 U292 ( .IN1(opA_EXE[13]), .IN2(n307), .IN3(n304), .IN4(fwd3[13]), 
        .IN5(n95), .Q(opA[13]) );
  AO22X1 U293 ( .IN1(fwd_opA[2]), .IN2(data_addr[13]), .IN3(n280), .IN4(
        reg_data_WB[13]), .Q(n95) );
  AO221X1 U294 ( .IN1(opA_EXE[12]), .IN2(n307), .IN3(n304), .IN4(fwd3[12]), 
        .IN5(n96), .Q(opA[12]) );
  AO22X1 U295 ( .IN1(fwd_opA[2]), .IN2(data_addr[12]), .IN3(n279), .IN4(
        reg_data_WB[12]), .Q(n96) );
  AO221X1 U296 ( .IN1(opA_EXE[11]), .IN2(n307), .IN3(n304), .IN4(fwd3[11]), 
        .IN5(n97), .Q(opA[11]) );
  AO22X1 U297 ( .IN1(fwd_opA[2]), .IN2(data_addr[11]), .IN3(n68), .IN4(
        reg_data_WB[11]), .Q(n97) );
  AO221X1 U298 ( .IN1(opA_EXE[10]), .IN2(n307), .IN3(n304), .IN4(fwd3[10]), 
        .IN5(n98), .Q(opA[10]) );
  AO22X1 U299 ( .IN1(fwd_opA[2]), .IN2(data_addr[10]), .IN3(n280), .IN4(
        reg_data_WB[10]), .Q(n98) );
  AO221X1 U300 ( .IN1(opA_EXE[0]), .IN2(n307), .IN3(n304), .IN4(fwd3[0]), 
        .IN5(n99), .Q(opA[0]) );
  AO22X1 U301 ( .IN1(fwd_opA[2]), .IN2(data_addr[0]), .IN3(n279), .IN4(
        reg_data_WB[0]), .Q(n99) );
  NAND4X0 U304 ( .IN1(n100), .IN2(n101), .IN3(n102), .IN4(n103), .QN(
        next_pc[9]) );
  AOI222X1 U305 ( .IN1(sel_pc[2]), .IN2(bra_pc[9]), .IN3(pc_p4_IF[9]), .IN4(
        n299), .IN5(n278), .IN6(imm_j[9]), .QN(n103) );
  AOI22X1 U306 ( .IN1(data_addr[9]), .IN2(n273), .IN3(reg_data_WB[9]), .IN4(
        n277), .QN(n102) );
  NAND4X0 U307 ( .IN1(n110), .IN2(n111), .IN3(n112), .IN4(n113), .QN(
        next_pc[8]) );
  AOI222X1 U308 ( .IN1(bra_pc[8]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[8]), .IN4(
        n301), .IN5(n105), .IN6(imm_alu[3]), .QN(n113) );
  AOI22X1 U309 ( .IN1(data_addr[8]), .IN2(n106), .IN3(reg_data_WB[8]), .IN4(
        n107), .QN(n112) );
  NAND4X0 U310 ( .IN1(n114), .IN2(n115), .IN3(n116), .IN4(n117), .QN(
        next_pc[7]) );
  AOI222X1 U311 ( .IN1(bra_pc[7]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[7]), .IN4(
        n301), .IN5(n278), .IN6(imm_alu[2]), .QN(n117) );
  AOI22X1 U312 ( .IN1(data_addr[7]), .IN2(n274), .IN3(reg_data_WB[7]), .IN4(
        n277), .QN(n116) );
  NAND4X0 U313 ( .IN1(n118), .IN2(n119), .IN3(n120), .IN4(n121), .QN(
        next_pc[6]) );
  AOI222X1 U314 ( .IN1(bra_pc[6]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[6]), .IN4(
        n301), .IN5(n105), .IN6(imm_alu[1]), .QN(n121) );
  AOI22X1 U315 ( .IN1(data_addr[6]), .IN2(n273), .IN3(reg_data_WB[6]), .IN4(
        n107), .QN(n120) );
  NAND4X0 U316 ( .IN1(n122), .IN2(n123), .IN3(n124), .IN4(n125), .QN(
        next_pc[5]) );
  AOI222X1 U317 ( .IN1(bra_pc[5]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[5]), .IN4(
        n301), .IN5(n278), .IN6(imm_alu[0]), .QN(n125) );
  AOI22X1 U318 ( .IN1(data_addr[5]), .IN2(n106), .IN3(reg_data_WB[5]), .IN4(
        n277), .QN(n124) );
  NAND4X0 U319 ( .IN1(n126), .IN2(n127), .IN3(n128), .IN4(n129), .QN(
        next_pc[4]) );
  AOI222X1 U320 ( .IN1(bra_pc[4]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[4]), .IN4(
        n301), .IN5(n105), .IN6(rd[4]), .QN(n129) );
  AOI22X1 U321 ( .IN1(data_addr[4]), .IN2(n274), .IN3(reg_data_WB[4]), .IN4(
        n107), .QN(n128) );
  NAND4X0 U322 ( .IN1(n130), .IN2(n131), .IN3(n132), .IN4(n133), .QN(
        next_pc[3]) );
  AOI222X1 U323 ( .IN1(bra_pc[3]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[3]), .IN4(
        n301), .IN5(n278), .IN6(rd[3]), .QN(n133) );
  AOI22X1 U324 ( .IN1(data_addr[3]), .IN2(n273), .IN3(reg_data_WB[3]), .IN4(
        n277), .QN(n132) );
  NAND4X0 U325 ( .IN1(n134), .IN2(n135), .IN3(n136), .IN4(n137), .QN(
        next_pc[31]) );
  AOI222X1 U326 ( .IN1(bra_pc[31]), .IN2(sel_pc[2]), .IN3(n107), .IN4(
        reg_data_WB[31]), .IN5(pc_p4_IF[31]), .IN6(n299), .QN(n137) );
  AOI22X1 U327 ( .IN1(fwd0[31]), .IN2(n295), .IN3(n274), .IN4(data_addr[31]), 
        .QN(n136) );
  NAND4X0 U328 ( .IN1(n138), .IN2(n135), .IN3(n139), .IN4(n140), .QN(
        next_pc[30]) );
  AOI222X1 U329 ( .IN1(bra_pc[30]), .IN2(sel_pc[2]), .IN3(n277), .IN4(
        reg_data_WB[30]), .IN5(pc_p4_IF[30]), .IN6(n299), .QN(n140) );
  AOI22X1 U330 ( .IN1(fwd0[30]), .IN2(n295), .IN3(n273), .IN4(data_addr[30]), 
        .QN(n139) );
  NAND4X0 U331 ( .IN1(n141), .IN2(n142), .IN3(n143), .IN4(n144), .QN(
        next_pc[2]) );
  AOI222X1 U332 ( .IN1(bra_pc[2]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[2]), .IN4(
        n300), .IN5(n105), .IN6(rd[2]), .QN(n144) );
  AOI22X1 U333 ( .IN1(data_addr[2]), .IN2(n106), .IN3(reg_data_WB[2]), .IN4(
        n107), .QN(n143) );
  NAND4X0 U334 ( .IN1(n145), .IN2(n135), .IN3(n146), .IN4(n147), .QN(
        next_pc[29]) );
  AOI222X1 U335 ( .IN1(bra_pc[29]), .IN2(sel_pc[2]), .IN3(n107), .IN4(
        reg_data_WB[29]), .IN5(pc_p4_IF[29]), .IN6(n299), .QN(n147) );
  AOI22X1 U336 ( .IN1(fwd0[29]), .IN2(n295), .IN3(n106), .IN4(data_addr[29]), 
        .QN(n146) );
  NAND4X0 U337 ( .IN1(n148), .IN2(n135), .IN3(n149), .IN4(n150), .QN(
        next_pc[28]) );
  AOI222X1 U338 ( .IN1(bra_pc[28]), .IN2(sel_pc[2]), .IN3(n277), .IN4(
        reg_data_WB[28]), .IN5(pc_p4_IF[28]), .IN6(n299), .QN(n150) );
  AOI22X1 U339 ( .IN1(fwd0[28]), .IN2(n295), .IN3(n274), .IN4(data_addr[28]), 
        .QN(n149) );
  NAND4X0 U340 ( .IN1(n151), .IN2(n135), .IN3(n152), .IN4(n153), .QN(
        next_pc[27]) );
  AOI222X1 U341 ( .IN1(bra_pc[27]), .IN2(sel_pc[2]), .IN3(n107), .IN4(
        reg_data_WB[27]), .IN5(pc_p4_IF[27]), .IN6(n299), .QN(n153) );
  AOI22X1 U342 ( .IN1(fwd0[27]), .IN2(n295), .IN3(n273), .IN4(data_addr[27]), 
        .QN(n152) );
  NAND4X0 U343 ( .IN1(n154), .IN2(n135), .IN3(n155), .IN4(n156), .QN(
        next_pc[26]) );
  AOI222X1 U344 ( .IN1(bra_pc[26]), .IN2(sel_pc[2]), .IN3(n277), .IN4(
        reg_data_WB[26]), .IN5(pc_p4_IF[26]), .IN6(n299), .QN(n156) );
  AOI22X1 U345 ( .IN1(fwd0[26]), .IN2(n295), .IN3(n106), .IN4(data_addr[26]), 
        .QN(n155) );
  NAND4X0 U346 ( .IN1(n157), .IN2(n135), .IN3(n158), .IN4(n159), .QN(
        next_pc[25]) );
  AOI222X1 U347 ( .IN1(bra_pc[25]), .IN2(sel_pc[2]), .IN3(n107), .IN4(
        reg_data_WB[25]), .IN5(pc_p4_IF[25]), .IN6(n299), .QN(n159) );
  AOI22X1 U348 ( .IN1(fwd0[25]), .IN2(n295), .IN3(n274), .IN4(data_addr[25]), 
        .QN(n158) );
  NAND4X0 U349 ( .IN1(n160), .IN2(n161), .IN3(n162), .IN4(n163), .QN(
        next_pc[24]) );
  AOI222X1 U350 ( .IN1(bra_pc[24]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[24]), .IN4(
        n300), .IN5(n278), .IN6(funct[5]), .QN(n163) );
  AOI22X1 U351 ( .IN1(data_addr[24]), .IN2(n274), .IN3(reg_data_WB[24]), .IN4(
        n277), .QN(n162) );
  NAND4X0 U352 ( .IN1(n164), .IN2(n165), .IN3(n166), .IN4(n167), .QN(
        next_pc[23]) );
  AOI222X1 U353 ( .IN1(bra_pc[23]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[23]), .IN4(
        n300), .IN5(n105), .IN6(funct[4]), .QN(n167) );
  AOI22X1 U354 ( .IN1(data_addr[23]), .IN2(n273), .IN3(reg_data_WB[23]), .IN4(
        n107), .QN(n166) );
  NAND4X0 U355 ( .IN1(n168), .IN2(n169), .IN3(n170), .IN4(n171), .QN(
        next_pc[22]) );
  AOI222X1 U356 ( .IN1(bra_pc[22]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[22]), .IN4(
        n300), .IN5(n278), .IN6(funct[3]), .QN(n171) );
  AOI22X1 U357 ( .IN1(data_addr[22]), .IN2(n106), .IN3(reg_data_WB[22]), .IN4(
        n277), .QN(n170) );
  NAND4X0 U358 ( .IN1(n172), .IN2(n173), .IN3(n174), .IN4(n175), .QN(
        next_pc[21]) );
  AOI222X1 U359 ( .IN1(bra_pc[21]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[21]), .IN4(
        n300), .IN5(n105), .IN6(funct[2]), .QN(n175) );
  AOI22X1 U360 ( .IN1(data_addr[21]), .IN2(n274), .IN3(reg_data_WB[21]), .IN4(
        n107), .QN(n174) );
  NAND4X0 U361 ( .IN1(n176), .IN2(n177), .IN3(n178), .IN4(n179), .QN(
        next_pc[20]) );
  AOI222X1 U362 ( .IN1(bra_pc[20]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[20]), .IN4(
        n300), .IN5(n278), .IN6(funct[1]), .QN(n179) );
  AOI22X1 U363 ( .IN1(data_addr[20]), .IN2(n273), .IN3(reg_data_WB[20]), .IN4(
        n277), .QN(n178) );
  NAND4X0 U364 ( .IN1(n180), .IN2(n181), .IN3(n182), .IN4(n183), .QN(
        next_pc[1]) );
  AOI222X1 U365 ( .IN1(bra_pc[1]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[1]), .IN4(
        n300), .IN5(n105), .IN6(rd[1]), .QN(n183) );
  AOI22X1 U366 ( .IN1(data_addr[1]), .IN2(n106), .IN3(reg_data_WB[1]), .IN4(
        n107), .QN(n182) );
  NAND4X0 U367 ( .IN1(n184), .IN2(n185), .IN3(n186), .IN4(n187), .QN(
        next_pc[19]) );
  AOI222X1 U368 ( .IN1(bra_pc[19]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[19]), .IN4(
        n300), .IN5(n278), .IN6(funct[0]), .QN(n187) );
  AOI22X1 U369 ( .IN1(data_addr[19]), .IN2(n274), .IN3(reg_data_WB[19]), .IN4(
        n277), .QN(n186) );
  NAND4X0 U370 ( .IN1(n188), .IN2(n189), .IN3(n190), .IN4(n191), .QN(
        next_pc[18]) );
  AOI222X1 U371 ( .IN1(bra_pc[18]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[18]), .IN4(
        n300), .IN5(n105), .IN6(imm_alu[8]), .QN(n191) );
  AOI22X1 U372 ( .IN1(data_addr[18]), .IN2(n273), .IN3(reg_data_WB[18]), .IN4(
        n107), .QN(n190) );
  NAND4X0 U373 ( .IN1(n192), .IN2(n193), .IN3(n194), .IN4(n195), .QN(
        next_pc[17]) );
  AOI222X1 U374 ( .IN1(bra_pc[17]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[17]), .IN4(
        n300), .IN5(n278), .IN6(imm_alu[7]), .QN(n195) );
  AOI22X1 U375 ( .IN1(data_addr[17]), .IN2(n106), .IN3(reg_data_WB[17]), .IN4(
        n277), .QN(n194) );
  NAND4X0 U376 ( .IN1(n196), .IN2(n197), .IN3(n198), .IN4(n199), .QN(
        next_pc[16]) );
  AOI222X1 U377 ( .IN1(bra_pc[16]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[16]), .IN4(
        n300), .IN5(n105), .IN6(imm_alu[6]), .QN(n199) );
  AOI22X1 U378 ( .IN1(data_addr[16]), .IN2(n274), .IN3(reg_data_WB[16]), .IN4(
        n107), .QN(n198) );
  NAND4X0 U379 ( .IN1(n200), .IN2(n201), .IN3(n202), .IN4(n203), .QN(
        next_pc[15]) );
  AOI222X1 U380 ( .IN1(bra_pc[15]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[15]), .IN4(
        n299), .IN5(n278), .IN6(imm_alu[5]), .QN(n203) );
  AOI22X1 U381 ( .IN1(data_addr[15]), .IN2(n273), .IN3(reg_data_WB[15]), .IN4(
        n277), .QN(n202) );
  NAND4X0 U382 ( .IN1(n204), .IN2(n205), .IN3(n206), .IN4(n207), .QN(
        next_pc[14]) );
  AOI222X1 U383 ( .IN1(bra_pc[14]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[14]), .IN4(
        n299), .IN5(n105), .IN6(imm_alu[4]), .QN(n207) );
  AOI22X1 U384 ( .IN1(data_addr[14]), .IN2(n106), .IN3(reg_data_WB[14]), .IN4(
        n107), .QN(n206) );
  NAND4X0 U385 ( .IN1(n208), .IN2(n209), .IN3(n210), .IN4(n211), .QN(
        next_pc[13]) );
  AOI222X1 U386 ( .IN1(bra_pc[13]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[13]), .IN4(
        n299), .IN5(n278), .IN6(imm_j[13]), .QN(n211) );
  AOI22X1 U387 ( .IN1(data_addr[13]), .IN2(n274), .IN3(reg_data_WB[13]), .IN4(
        n277), .QN(n210) );
  NAND4X0 U388 ( .IN1(n212), .IN2(n213), .IN3(n214), .IN4(n215), .QN(
        next_pc[12]) );
  AOI222X1 U389 ( .IN1(bra_pc[12]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[12]), .IN4(
        n299), .IN5(n105), .IN6(imm_j[12]), .QN(n215) );
  AOI22X1 U390 ( .IN1(data_addr[12]), .IN2(n273), .IN3(reg_data_WB[12]), .IN4(
        n107), .QN(n214) );
  NAND4X0 U391 ( .IN1(n216), .IN2(n217), .IN3(n218), .IN4(n219), .QN(
        next_pc[11]) );
  AOI222X1 U392 ( .IN1(bra_pc[11]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[11]), .IN4(
        n300), .IN5(n278), .IN6(imm_j[11]), .QN(n219) );
  AOI22X1 U393 ( .IN1(data_addr[11]), .IN2(n106), .IN3(reg_data_WB[11]), .IN4(
        n277), .QN(n218) );
  NAND4X0 U394 ( .IN1(n220), .IN2(n221), .IN3(n222), .IN4(n223), .QN(
        next_pc[10]) );
  AOI222X1 U395 ( .IN1(bra_pc[10]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[10]), .IN4(
        n299), .IN5(n105), .IN6(imm_j[10]), .QN(n223) );
  AOI22X1 U396 ( .IN1(data_addr[10]), .IN2(n274), .IN3(reg_data_WB[10]), .IN4(
        n107), .QN(n222) );
  NAND4X0 U397 ( .IN1(n224), .IN2(n225), .IN3(n226), .IN4(n227), .QN(
        next_pc[0]) );
  AOI222X1 U398 ( .IN1(bra_pc[0]), .IN2(sel_pc[2]), .IN3(pc_p4_IF[0]), .IN4(
        n300), .IN5(n278), .IN6(rd[0]), .QN(n227) );
  AOI22X1 U400 ( .IN1(data_addr[0]), .IN2(n273), .IN3(reg_data_WB[0]), .IN4(
        n277), .QN(n226) );
  AND3X1 U401 ( .IN1(n318), .IN2(n321), .IN3(fwd_jr[1]), .Q(n106) );
  NAND3X0 U404 ( .IN1(n323), .IN2(n317), .IN3(sel_pc[0]), .QN(n228) );
  AO221X1 U405 ( .IN1(mem_data_EXE0[9]), .IN2(n290), .IN3(n287), .IN4(fwd3[9]), 
        .IN5(n231), .Q(mem_data_EXE[9]) );
  AO22X1 U406 ( .IN1(fwd_sw[2]), .IN2(data_addr[9]), .IN3(n276), .IN4(
        reg_data_WB[9]), .Q(n231) );
  AO221X1 U407 ( .IN1(mem_data_EXE0[8]), .IN2(n290), .IN3(n287), .IN4(fwd3[8]), 
        .IN5(n233), .Q(mem_data_EXE[8]) );
  AO22X1 U408 ( .IN1(fwd_sw[2]), .IN2(data_addr[8]), .IN3(n275), .IN4(
        reg_data_WB[8]), .Q(n233) );
  AO221X1 U409 ( .IN1(mem_data_EXE0[7]), .IN2(n290), .IN3(n287), .IN4(fwd3[7]), 
        .IN5(n234), .Q(mem_data_EXE[7]) );
  AO22X1 U410 ( .IN1(fwd_sw[2]), .IN2(data_addr[7]), .IN3(n232), .IN4(
        reg_data_WB[7]), .Q(n234) );
  AO221X1 U411 ( .IN1(mem_data_EXE0[6]), .IN2(n290), .IN3(n287), .IN4(fwd3[6]), 
        .IN5(n235), .Q(mem_data_EXE[6]) );
  AO22X1 U412 ( .IN1(fwd_sw[2]), .IN2(data_addr[6]), .IN3(n276), .IN4(
        reg_data_WB[6]), .Q(n235) );
  AO221X1 U413 ( .IN1(mem_data_EXE0[5]), .IN2(n290), .IN3(n287), .IN4(fwd3[5]), 
        .IN5(n236), .Q(mem_data_EXE[5]) );
  AO22X1 U414 ( .IN1(fwd_sw[2]), .IN2(data_addr[5]), .IN3(n275), .IN4(
        reg_data_WB[5]), .Q(n236) );
  AO221X1 U415 ( .IN1(mem_data_EXE0[4]), .IN2(n290), .IN3(n287), .IN4(fwd3[4]), 
        .IN5(n237), .Q(mem_data_EXE[4]) );
  AO22X1 U416 ( .IN1(fwd_sw[2]), .IN2(data_addr[4]), .IN3(n232), .IN4(
        reg_data_WB[4]), .Q(n237) );
  AO221X1 U417 ( .IN1(mem_data_EXE0[3]), .IN2(n290), .IN3(n287), .IN4(fwd3[3]), 
        .IN5(n238), .Q(mem_data_EXE[3]) );
  AO22X1 U418 ( .IN1(fwd_sw[2]), .IN2(data_addr[3]), .IN3(n276), .IN4(
        reg_data_WB[3]), .Q(n238) );
  AO221X1 U419 ( .IN1(mem_data_EXE0[31]), .IN2(n290), .IN3(n287), .IN4(
        fwd3[31]), .IN5(n239), .Q(mem_data_EXE[31]) );
  AO22X1 U420 ( .IN1(fwd_sw[2]), .IN2(data_addr[31]), .IN3(n275), .IN4(
        reg_data_WB[31]), .Q(n239) );
  AO221X1 U421 ( .IN1(mem_data_EXE0[30]), .IN2(n290), .IN3(n287), .IN4(
        fwd3[30]), .IN5(n240), .Q(mem_data_EXE[30]) );
  AO22X1 U422 ( .IN1(fwd_sw[2]), .IN2(data_addr[30]), .IN3(n232), .IN4(
        reg_data_WB[30]), .Q(n240) );
  AO221X1 U423 ( .IN1(mem_data_EXE0[2]), .IN2(n290), .IN3(n287), .IN4(fwd3[2]), 
        .IN5(n241), .Q(mem_data_EXE[2]) );
  AO22X1 U424 ( .IN1(fwd_sw[2]), .IN2(data_addr[2]), .IN3(n276), .IN4(
        reg_data_WB[2]), .Q(n241) );
  AO221X1 U425 ( .IN1(mem_data_EXE0[29]), .IN2(n290), .IN3(n287), .IN4(
        fwd3[29]), .IN5(n242), .Q(mem_data_EXE[29]) );
  AO22X1 U426 ( .IN1(fwd_sw[2]), .IN2(data_addr[29]), .IN3(n275), .IN4(
        reg_data_WB[29]), .Q(n242) );
  AO221X1 U427 ( .IN1(mem_data_EXE0[28]), .IN2(n290), .IN3(n287), .IN4(
        fwd3[28]), .IN5(n243), .Q(mem_data_EXE[28]) );
  AO22X1 U428 ( .IN1(fwd_sw[2]), .IN2(data_addr[28]), .IN3(n232), .IN4(
        reg_data_WB[28]), .Q(n243) );
  AO221X1 U429 ( .IN1(mem_data_EXE0[27]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[27]), .IN5(n244), .Q(mem_data_EXE[27]) );
  AO22X1 U430 ( .IN1(fwd_sw[2]), .IN2(data_addr[27]), .IN3(n276), .IN4(
        reg_data_WB[27]), .Q(n244) );
  AO221X1 U431 ( .IN1(mem_data_EXE0[26]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[26]), .IN5(n245), .Q(mem_data_EXE[26]) );
  AO22X1 U432 ( .IN1(fwd_sw[2]), .IN2(data_addr[26]), .IN3(n275), .IN4(
        reg_data_WB[26]), .Q(n245) );
  AO221X1 U433 ( .IN1(mem_data_EXE0[25]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[25]), .IN5(n246), .Q(mem_data_EXE[25]) );
  AO22X1 U434 ( .IN1(fwd_sw[2]), .IN2(data_addr[25]), .IN3(n232), .IN4(
        reg_data_WB[25]), .Q(n246) );
  AO221X1 U435 ( .IN1(mem_data_EXE0[24]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[24]), .IN5(n247), .Q(mem_data_EXE[24]) );
  AO22X1 U436 ( .IN1(fwd_sw[2]), .IN2(data_addr[24]), .IN3(n276), .IN4(
        reg_data_WB[24]), .Q(n247) );
  AO221X1 U437 ( .IN1(mem_data_EXE0[23]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[23]), .IN5(n248), .Q(mem_data_EXE[23]) );
  AO22X1 U438 ( .IN1(fwd_sw[2]), .IN2(data_addr[23]), .IN3(n275), .IN4(
        reg_data_WB[23]), .Q(n248) );
  AO221X1 U439 ( .IN1(mem_data_EXE0[22]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[22]), .IN5(n249), .Q(mem_data_EXE[22]) );
  AO22X1 U440 ( .IN1(fwd_sw[2]), .IN2(data_addr[22]), .IN3(n232), .IN4(
        reg_data_WB[22]), .Q(n249) );
  AO221X1 U441 ( .IN1(mem_data_EXE0[21]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[21]), .IN5(n250), .Q(mem_data_EXE[21]) );
  AO22X1 U442 ( .IN1(fwd_sw[2]), .IN2(data_addr[21]), .IN3(n276), .IN4(
        reg_data_WB[21]), .Q(n250) );
  AO221X1 U443 ( .IN1(mem_data_EXE0[20]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[20]), .IN5(n251), .Q(mem_data_EXE[20]) );
  AO22X1 U444 ( .IN1(fwd_sw[2]), .IN2(data_addr[20]), .IN3(n275), .IN4(
        reg_data_WB[20]), .Q(n251) );
  AO221X1 U445 ( .IN1(mem_data_EXE0[1]), .IN2(n291), .IN3(n288), .IN4(fwd3[1]), 
        .IN5(n252), .Q(mem_data_EXE[1]) );
  AO22X1 U446 ( .IN1(fwd_sw[2]), .IN2(data_addr[1]), .IN3(n232), .IN4(
        reg_data_WB[1]), .Q(n252) );
  AO221X1 U447 ( .IN1(mem_data_EXE0[19]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[19]), .IN5(n253), .Q(mem_data_EXE[19]) );
  AO22X1 U448 ( .IN1(fwd_sw[2]), .IN2(data_addr[19]), .IN3(n276), .IN4(
        reg_data_WB[19]), .Q(n253) );
  AO221X1 U449 ( .IN1(mem_data_EXE0[18]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[18]), .IN5(n254), .Q(mem_data_EXE[18]) );
  AO22X1 U450 ( .IN1(fwd_sw[2]), .IN2(data_addr[18]), .IN3(n275), .IN4(
        reg_data_WB[18]), .Q(n254) );
  AO221X1 U451 ( .IN1(mem_data_EXE0[17]), .IN2(n291), .IN3(n288), .IN4(
        fwd3[17]), .IN5(n255), .Q(mem_data_EXE[17]) );
  AO22X1 U452 ( .IN1(fwd_sw[2]), .IN2(data_addr[17]), .IN3(n232), .IN4(
        reg_data_WB[17]), .Q(n255) );
  AO221X1 U453 ( .IN1(mem_data_EXE0[16]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[16]), .IN5(n256), .Q(mem_data_EXE[16]) );
  AO22X1 U454 ( .IN1(fwd_sw[2]), .IN2(data_addr[16]), .IN3(n276), .IN4(
        reg_data_WB[16]), .Q(n256) );
  AO221X1 U455 ( .IN1(mem_data_EXE0[15]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[15]), .IN5(n257), .Q(mem_data_EXE[15]) );
  AO22X1 U456 ( .IN1(fwd_sw[2]), .IN2(data_addr[15]), .IN3(n275), .IN4(
        reg_data_WB[15]), .Q(n257) );
  AO221X1 U457 ( .IN1(mem_data_EXE0[14]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[14]), .IN5(n258), .Q(mem_data_EXE[14]) );
  AO22X1 U458 ( .IN1(fwd_sw[2]), .IN2(data_addr[14]), .IN3(n232), .IN4(
        reg_data_WB[14]), .Q(n258) );
  AO221X1 U459 ( .IN1(mem_data_EXE0[13]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[13]), .IN5(n259), .Q(mem_data_EXE[13]) );
  AO22X1 U460 ( .IN1(fwd_sw[2]), .IN2(data_addr[13]), .IN3(n276), .IN4(
        reg_data_WB[13]), .Q(n259) );
  AO221X1 U461 ( .IN1(mem_data_EXE0[12]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[12]), .IN5(n260), .Q(mem_data_EXE[12]) );
  AO22X1 U462 ( .IN1(fwd_sw[2]), .IN2(data_addr[12]), .IN3(n275), .IN4(
        reg_data_WB[12]), .Q(n260) );
  AO221X1 U463 ( .IN1(mem_data_EXE0[11]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[11]), .IN5(n261), .Q(mem_data_EXE[11]) );
  AO22X1 U464 ( .IN1(fwd_sw[2]), .IN2(data_addr[11]), .IN3(n232), .IN4(
        reg_data_WB[11]), .Q(n261) );
  AO221X1 U465 ( .IN1(mem_data_EXE0[10]), .IN2(n292), .IN3(n289), .IN4(
        fwd3[10]), .IN5(n262), .Q(mem_data_EXE[10]) );
  AO22X1 U466 ( .IN1(fwd_sw[2]), .IN2(data_addr[10]), .IN3(n276), .IN4(
        reg_data_WB[10]), .Q(n262) );
  AO221X1 U467 ( .IN1(mem_data_EXE0[0]), .IN2(n292), .IN3(n289), .IN4(fwd3[0]), 
        .IN5(n263), .Q(mem_data_EXE[0]) );
  AO22X1 U468 ( .IN1(fwd_sw[2]), .IN2(data_addr[0]), .IN3(n275), .IN4(
        reg_data_WB[0]), .Q(n263) );
  reg32_0 PC ( .clk(clk), .nrst(nrst), .en(n319), .data_in(next_pc), 
        .data_out(pc_IF) );
  if_id_reg IF_ID ( .clk(clk), .nrst(nrst), .en(n319), .flush(flush[1]), 
        .cur_pc0(pc_IF), .next_pc0(pc_p4_IF), .cur_pc(pc_ID), .next_pc(
        pc_p4_ID) );
  rf RF ( .clk(clk), .nrst(nrst), .wr_en(wr_rf), .rd_addrA(rs1), .rd_addrB(rs2), .wr_addr(reg_addr_WB), .wr_data(reg_data_WB), .rd_dataA(opA_ID), .rd_dataB(
        mem_data_ID) );
  id_exe_reg ID_EXE ( .clk(clk), .nrst(nrst), .en(n319), .flush(flush[0]), 
        .cur_pc0(pc_ID), .next_pc0(pc_p4_ID), .bra_off0({funct[6], funct[6], 
        funct[6], funct[6], funct[6], funct[6], funct[6], funct[6], funct[6], 
        funct[6], funct[6], funct[6], funct[6], funct[6], funct[6], funct[6], 
        funct, imm_alu[3:0], rd}), .opA0(opA_ID), .opB0(opB_ID), .mem_data0(
        mem_data_ID), .reg_addr0(reg_addr_ID), .cur_pc(pc_EXE), .next_pc(
        pc_p4_EXE), .bra_off(bra_off_EXE), .opA(opA_EXE), .opB(opB_EXE), 
        .mem_data(mem_data_EXE0), .reg_addr(reg_addr_EXE) );
  alu ALU ( .opA(opA), .opB(opB), .res(fwd0), .alu_code(alu_code), .z(zero) );
  exe_mem_reg EXE_MEM ( .clk(clk), .nrst(nrst), .cur_pc0(pc_EXE), .next_pc0(
        pc_p4_EXE), .alu_out0(fwd0), .mem_data0(mem_data_EXE), .reg_addr0(
        reg_addr_EXE), .cur_pc(pc_MEM), .next_pc(pc_p4_MEM), .alu_out(
        data_addr), .mem_data(data_out), .reg_addr(reg_addr_MEM) );
  mem_wb_reg MEM_WB ( .clk(clk), .nrst(nrst), .cur_pc0(pc_MEM), .next_pc0(
        pc_p4_MEM), .reg_data0(reg_data_MEM), .reg_addr0(reg_addr_MEM), 
        .cur_pc(pc_WB), .reg_data(reg_data_WB), .reg_addr(reg_addr_WB) );
  reg32_5 FWD_WB ( .clk(clk), .nrst(nrst), .en(1'b1), .data_in(reg_data_WB), 
        .data_out(fwd3) );
  control CTRL ( .clk(clk), .nrst(nrst), .zero(zero), .inst(inst), .jr(jr), 
        .jal(jal), .jal_pc(jal_pc), .load(load), .wr_mem(data_wr), .use_imm(
        use_imm), .sw(sw), .debug_inst({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, funct, imm_alu[8:4], imm_j, imm_alu[3:0], rd, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133}), .alu_code(
        alu_code), .sel_pc(sel_pc), .flush(flush), .wr_rf(wr_rf), .stall(stall), .fwd_opA(fwd_opA), .fwd_opB(fwd_opB), .fwd_sw(fwd_sw), .fwd_jr(fwd_jr) );
  pipeline_riscv_DW01_add_0 add_151 ( .A(pc_p4_EXE), .B(bra_off_EXE), .CI(1'b0), .SUM(bra_pc) );
  pipeline_riscv_DW01_add_1 add_76 ( .A(pc_IF), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_p4_IF) );
  OR3X1 U471 ( .IN1(sel_pc[1]), .IN2(sel_pc[2]), .IN3(sel_pc[0]), .Q(n264) );
  OR3X1 U472 ( .IN1(fwd_opA[1]), .IN2(fwd_opA[2]), .IN3(n330), .Q(n265) );
  OR3X1 U473 ( .IN1(fwd_opA[1]), .IN2(fwd_opA[2]), .IN3(fwd_opA[0]), .Q(n266)
         );
  OR3X1 U474 ( .IN1(fwd_opB[1]), .IN2(fwd_opB[2]), .IN3(n326), .Q(n267) );
  OR3X1 U475 ( .IN1(fwd_opB[1]), .IN2(fwd_opB[2]), .IN3(fwd_opB[0]), .Q(n268)
         );
  OR4X1 U476 ( .IN1(n228), .IN2(fwd_jr[0]), .IN3(fwd_jr[1]), .IN4(fwd_jr[2]), 
        .Q(n269) );
  OR4X1 U477 ( .IN1(n320), .IN2(n228), .IN3(fwd_jr[1]), .IN4(fwd_jr[2]), .Q(
        n270) );
  OR3X1 U478 ( .IN1(fwd_sw[1]), .IN2(fwd_sw[2]), .IN3(n328), .Q(n271) );
  OR3X1 U479 ( .IN1(fwd_sw[1]), .IN2(fwd_sw[2]), .IN3(fwd_sw[0]), .Q(n272) );
  INVX0 U480 ( .INP(sel_pc[2]), .ZN(n317) );
  INVX0 U481 ( .INP(jal), .ZN(n316) );
  INVX0 U482 ( .INP(n269), .ZN(n298) );
  INVX0 U483 ( .INP(n270), .ZN(n295) );
  NAND2X1 U484 ( .IN1(fwd0[9]), .IN2(n295), .QN(n100) );
  INVX0 U485 ( .INP(n270), .ZN(n293) );
  INVX0 U486 ( .INP(n270), .ZN(n294) );
  INVX0 U487 ( .INP(n269), .ZN(n296) );
  INVX0 U488 ( .INP(n269), .ZN(n297) );
  NAND2X1 U489 ( .IN1(fwd0[1]), .IN2(n293), .QN(n180) );
  NAND2X1 U490 ( .IN1(fwd0[12]), .IN2(n293), .QN(n212) );
  NAND2X1 U491 ( .IN1(fwd0[16]), .IN2(n293), .QN(n196) );
  NAND2X1 U492 ( .IN1(fwd0[23]), .IN2(n294), .QN(n164) );
  NAND2X1 U493 ( .IN1(fwd0[10]), .IN2(n293), .QN(n220) );
  NAND2X1 U494 ( .IN1(fwd0[14]), .IN2(n293), .QN(n204) );
  NAND2X1 U495 ( .IN1(fwd0[18]), .IN2(n293), .QN(n188) );
  NAND2X1 U496 ( .IN1(fwd0[21]), .IN2(n294), .QN(n172) );
  NAND2X1 U497 ( .IN1(fwd0[13]), .IN2(n293), .QN(n208) );
  NAND2X1 U498 ( .IN1(fwd0[17]), .IN2(n293), .QN(n192) );
  NAND2X1 U499 ( .IN1(fwd0[20]), .IN2(n294), .QN(n176) );
  NAND2X1 U500 ( .IN1(fwd0[24]), .IN2(n294), .QN(n160) );
  NAND2X1 U501 ( .IN1(fwd0[2]), .IN2(n294), .QN(n141) );
  NAND2X1 U502 ( .IN1(fwd0[11]), .IN2(n293), .QN(n216) );
  NAND2X1 U503 ( .IN1(fwd0[15]), .IN2(n293), .QN(n200) );
  NAND2X1 U504 ( .IN1(fwd0[19]), .IN2(n293), .QN(n184) );
  NAND2X1 U505 ( .IN1(fwd0[22]), .IN2(n294), .QN(n168) );
  NOR2X0 U506 ( .IN1(n323), .IN2(sel_pc[2]), .QN(n105) );
  NOR2X0 U507 ( .IN1(n323), .IN2(sel_pc[2]), .QN(n278) );
  INVX0 U508 ( .INP(fwd_jr[0]), .ZN(n320) );
  INVX0 U509 ( .INP(n264), .ZN(n301) );
  INVX0 U510 ( .INP(n228), .ZN(n318) );
  NAND2X1 U511 ( .IN1(fwd0[0]), .IN2(n293), .QN(n224) );
  INVX0 U512 ( .INP(n264), .ZN(n299) );
  INVX0 U513 ( .INP(n264), .ZN(n300) );
  NOR2X0 U514 ( .IN1(n321), .IN2(n228), .QN(n107) );
  NOR2X0 U515 ( .IN1(n321), .IN2(n228), .QN(n277) );
  INVX0 U516 ( .INP(sel_pc[1]), .ZN(n323) );
  INVX0 U517 ( .INP(fwd_jr[2]), .ZN(n321) );
  INVX0 U518 ( .INP(n24), .ZN(n322) );
  INVX0 U519 ( .INP(jal_pc), .ZN(n324) );
  INVX0 U520 ( .INP(n316), .ZN(n315) );
  INVX0 U521 ( .INP(n316), .ZN(n314) );
  INVX0 U522 ( .INP(n267), .ZN(n310) );
  INVX0 U523 ( .INP(n265), .ZN(n304) );
  INVX0 U524 ( .INP(n268), .ZN(n313) );
  INVX0 U525 ( .INP(n266), .ZN(n307) );
  NAND2X1 U526 ( .IN1(n298), .IN2(mem_data_ID[3]), .QN(n131) );
  NAND2X1 U527 ( .IN1(n298), .IN2(mem_data_ID[4]), .QN(n127) );
  NAND2X1 U528 ( .IN1(n298), .IN2(mem_data_ID[5]), .QN(n123) );
  NAND2X1 U529 ( .IN1(n298), .IN2(mem_data_ID[6]), .QN(n119) );
  NAND2X1 U530 ( .IN1(n298), .IN2(mem_data_ID[7]), .QN(n115) );
  NAND2X1 U531 ( .IN1(n298), .IN2(mem_data_ID[8]), .QN(n111) );
  NAND2X1 U532 ( .IN1(n298), .IN2(mem_data_ID[9]), .QN(n101) );
  INVX0 U533 ( .INP(n267), .ZN(n309) );
  INVX0 U534 ( .INP(n267), .ZN(n308) );
  INVX0 U535 ( .INP(n265), .ZN(n303) );
  INVX0 U536 ( .INP(n265), .ZN(n302) );
  INVX0 U537 ( .INP(n268), .ZN(n312) );
  INVX0 U538 ( .INP(n266), .ZN(n306) );
  INVX0 U539 ( .INP(n268), .ZN(n311) );
  INVX0 U540 ( .INP(n266), .ZN(n305) );
  NOR2X0 U541 ( .IN1(jr), .IN2(sw), .QN(n24) );
  INVX0 U542 ( .INP(stall), .ZN(n319) );
  NOR2X0 U543 ( .IN1(n324), .IN2(load), .QN(n25) );
  NOR2X0 U544 ( .IN1(n324), .IN2(load), .QN(n284) );
  NOR2X0 U545 ( .IN1(jal_pc), .IN2(load), .QN(n286) );
  NOR2X0 U546 ( .IN1(jal_pc), .IN2(load), .QN(n285) );
  NOR2X0 U547 ( .IN1(jal_pc), .IN2(load), .QN(n26) );
  NOR2X0 U548 ( .IN1(n314), .IN2(use_imm), .QN(n28) );
  NOR2X0 U549 ( .IN1(n314), .IN2(use_imm), .QN(n283) );
  AND2X1 U550 ( .IN1(use_imm), .IN2(n316), .Q(n27) );
  INVX0 U551 ( .INP(n271), .ZN(n289) );
  INVX0 U552 ( .INP(n272), .ZN(n292) );
  INVX0 U553 ( .INP(n271), .ZN(n288) );
  INVX0 U554 ( .INP(n271), .ZN(n287) );
  INVX0 U555 ( .INP(n272), .ZN(n291) );
  INVX0 U556 ( .INP(n272), .ZN(n290) );
  NOR2X0 U557 ( .IN1(n325), .IN2(fwd_opB[2]), .QN(n281) );
  INVX0 U558 ( .INP(fwd_opB[0]), .ZN(n326) );
  INVX0 U559 ( .INP(fwd_opA[0]), .ZN(n330) );
  NAND2X1 U560 ( .IN1(n297), .IN2(mem_data_ID[25]), .QN(n157) );
  NAND2X1 U561 ( .IN1(n297), .IN2(mem_data_ID[26]), .QN(n154) );
  NAND2X1 U562 ( .IN1(n297), .IN2(mem_data_ID[27]), .QN(n151) );
  NAND2X1 U563 ( .IN1(n297), .IN2(mem_data_ID[28]), .QN(n148) );
  NAND2X1 U564 ( .IN1(n297), .IN2(mem_data_ID[29]), .QN(n145) );
  NAND2X1 U565 ( .IN1(n297), .IN2(mem_data_ID[30]), .QN(n138) );
  NAND2X1 U566 ( .IN1(n298), .IN2(mem_data_ID[31]), .QN(n134) );
  NAND2X1 U567 ( .IN1(n296), .IN2(mem_data_ID[0]), .QN(n225) );
  NAND2X1 U568 ( .IN1(n296), .IN2(mem_data_ID[1]), .QN(n181) );
  NAND2X1 U569 ( .IN1(n297), .IN2(mem_data_ID[2]), .QN(n142) );
  NAND2X1 U570 ( .IN1(fwd0[3]), .IN2(n294), .QN(n130) );
  NAND2X1 U571 ( .IN1(fwd0[4]), .IN2(n294), .QN(n126) );
  NAND2X1 U572 ( .IN1(fwd0[5]), .IN2(n294), .QN(n122) );
  NAND2X1 U573 ( .IN1(fwd0[6]), .IN2(n294), .QN(n118) );
  NAND2X1 U574 ( .IN1(fwd0[7]), .IN2(n294), .QN(n114) );
  NAND2X1 U575 ( .IN1(fwd0[8]), .IN2(n294), .QN(n110) );
  NAND2X1 U576 ( .IN1(n296), .IN2(mem_data_ID[10]), .QN(n221) );
  NAND2X1 U577 ( .IN1(n296), .IN2(mem_data_ID[11]), .QN(n217) );
  NAND2X1 U578 ( .IN1(n296), .IN2(mem_data_ID[12]), .QN(n213) );
  NAND2X1 U579 ( .IN1(n296), .IN2(mem_data_ID[13]), .QN(n209) );
  NAND2X1 U580 ( .IN1(n296), .IN2(mem_data_ID[14]), .QN(n205) );
  NAND2X1 U581 ( .IN1(n296), .IN2(mem_data_ID[15]), .QN(n201) );
  NAND2X1 U582 ( .IN1(n296), .IN2(mem_data_ID[16]), .QN(n197) );
  NAND2X1 U583 ( .IN1(n296), .IN2(mem_data_ID[17]), .QN(n193) );
  NAND2X1 U584 ( .IN1(n296), .IN2(mem_data_ID[18]), .QN(n189) );
  NAND2X1 U585 ( .IN1(n296), .IN2(mem_data_ID[19]), .QN(n185) );
  NAND2X1 U586 ( .IN1(n297), .IN2(mem_data_ID[20]), .QN(n177) );
  NAND2X1 U587 ( .IN1(n297), .IN2(mem_data_ID[21]), .QN(n173) );
  NAND2X1 U588 ( .IN1(n297), .IN2(mem_data_ID[22]), .QN(n169) );
  NAND2X1 U589 ( .IN1(n297), .IN2(mem_data_ID[23]), .QN(n165) );
  NAND2X1 U590 ( .IN1(n297), .IN2(mem_data_ID[24]), .QN(n161) );
  NOR2X0 U591 ( .IN1(n325), .IN2(fwd_opB[2]), .QN(n282) );
  NOR2X0 U592 ( .IN1(n329), .IN2(fwd_opA[2]), .QN(n279) );
  NOR2X0 U593 ( .IN1(n329), .IN2(fwd_opA[2]), .QN(n280) );
  NOR2X0 U594 ( .IN1(n325), .IN2(fwd_opB[2]), .QN(n33) );
  NOR2X0 U595 ( .IN1(n329), .IN2(fwd_opA[2]), .QN(n68) );
  NAND2X1 U596 ( .IN1(n105), .IN2(funct[6]), .QN(n135) );
  INVX0 U597 ( .INP(fwd_opB[1]), .ZN(n325) );
  INVX0 U598 ( .INP(fwd_opA[1]), .ZN(n329) );
  NOR2X0 U599 ( .IN1(n327), .IN2(fwd_sw[2]), .QN(n276) );
  NOR2X0 U600 ( .IN1(n327), .IN2(fwd_sw[2]), .QN(n275) );
  NOR2X0 U601 ( .IN1(n327), .IN2(fwd_sw[2]), .QN(n232) );
  AND2X1 U602 ( .IN1(funct[6]), .IN2(n27), .Q(n29) );
  INVX0 U603 ( .INP(fwd_sw[0]), .ZN(n328) );
  INVX0 U604 ( .INP(fwd_sw[1]), .ZN(n327) );
  AND3X1 U605 ( .IN1(n318), .IN2(n321), .IN3(fwd_jr[1]), .Q(n273) );
  AND3X1 U606 ( .IN1(n318), .IN2(n321), .IN3(fwd_jr[1]), .Q(n274) );
endmodule

